-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity fill_input is -- 
  generic (tag_length : integer); 
  port ( -- 
    system_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    system_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    system_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    writeModule1_call_reqs : out  std_logic_vector(0 downto 0);
    writeModule1_call_acks : in   std_logic_vector(0 downto 0);
    writeModule1_call_data : out  std_logic_vector(95 downto 0);
    writeModule1_call_tag  :  out  std_logic_vector(0 downto 0);
    writeModule1_return_reqs : out  std_logic_vector(0 downto 0);
    writeModule1_return_acks : in   std_logic_vector(0 downto 0);
    writeModule1_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity fill_input;
architecture fill_input_arch of fill_input is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal fill_input_CP_122_start: Boolean;
  signal fill_input_CP_122_symbol: Boolean;
  -- volatile/operator module components. 
  component writeModule1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      address : in  std_logic_vector(31 downto 0);
      data : in  std_logic_vector(63 downto 0);
      memoryModule_call_reqs : out  std_logic_vector(0 downto 0);
      memoryModule_call_acks : in   std_logic_vector(0 downto 0);
      memoryModule_call_data : out  std_logic_vector(96 downto 0);
      memoryModule_call_tag  :  out  std_logic_vector(0 downto 0);
      memoryModule_return_reqs : out  std_logic_vector(0 downto 0);
      memoryModule_return_acks : in   std_logic_vector(0 downto 0);
      memoryModule_return_data : in   std_logic_vector(63 downto 0);
      memoryModule_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal type_cast_138_inst_req_0 : boolean;
  signal type_cast_138_inst_ack_0 : boolean;
  signal type_cast_138_inst_req_1 : boolean;
  signal type_cast_138_inst_ack_1 : boolean;
  signal RPIPE_system_input_pipe_85_inst_req_0 : boolean;
  signal RPIPE_system_input_pipe_85_inst_ack_0 : boolean;
  signal RPIPE_system_input_pipe_85_inst_req_1 : boolean;
  signal RPIPE_system_input_pipe_85_inst_ack_1 : boolean;
  signal type_cast_89_inst_req_0 : boolean;
  signal type_cast_89_inst_ack_0 : boolean;
  signal type_cast_89_inst_req_1 : boolean;
  signal type_cast_89_inst_ack_1 : boolean;
  signal RPIPE_system_input_pipe_98_inst_req_0 : boolean;
  signal RPIPE_system_input_pipe_98_inst_ack_0 : boolean;
  signal RPIPE_system_input_pipe_98_inst_req_1 : boolean;
  signal RPIPE_system_input_pipe_98_inst_ack_1 : boolean;
  signal type_cast_102_inst_req_0 : boolean;
  signal type_cast_102_inst_ack_0 : boolean;
  signal type_cast_102_inst_req_1 : boolean;
  signal type_cast_102_inst_ack_1 : boolean;
  signal RPIPE_system_input_pipe_116_inst_req_0 : boolean;
  signal RPIPE_system_input_pipe_116_inst_ack_0 : boolean;
  signal RPIPE_system_input_pipe_116_inst_req_1 : boolean;
  signal RPIPE_system_input_pipe_116_inst_ack_1 : boolean;
  signal type_cast_120_inst_req_0 : boolean;
  signal type_cast_120_inst_ack_0 : boolean;
  signal type_cast_120_inst_req_1 : boolean;
  signal type_cast_120_inst_ack_1 : boolean;
  signal RPIPE_system_input_pipe_134_inst_req_0 : boolean;
  signal RPIPE_system_input_pipe_134_inst_ack_0 : boolean;
  signal RPIPE_system_input_pipe_134_inst_req_1 : boolean;
  signal RPIPE_system_input_pipe_134_inst_ack_1 : boolean;
  signal RPIPE_system_input_pipe_152_inst_req_0 : boolean;
  signal RPIPE_system_input_pipe_152_inst_ack_0 : boolean;
  signal RPIPE_system_input_pipe_152_inst_req_1 : boolean;
  signal RPIPE_system_input_pipe_152_inst_ack_1 : boolean;
  signal type_cast_156_inst_req_0 : boolean;
  signal type_cast_156_inst_ack_0 : boolean;
  signal type_cast_156_inst_req_1 : boolean;
  signal type_cast_156_inst_ack_1 : boolean;
  signal RPIPE_system_input_pipe_170_inst_req_0 : boolean;
  signal RPIPE_system_input_pipe_170_inst_ack_0 : boolean;
  signal RPIPE_system_input_pipe_170_inst_req_1 : boolean;
  signal RPIPE_system_input_pipe_170_inst_ack_1 : boolean;
  signal type_cast_174_inst_req_0 : boolean;
  signal type_cast_174_inst_ack_0 : boolean;
  signal type_cast_174_inst_req_1 : boolean;
  signal type_cast_174_inst_ack_1 : boolean;
  signal RPIPE_system_input_pipe_188_inst_req_0 : boolean;
  signal RPIPE_system_input_pipe_188_inst_ack_0 : boolean;
  signal RPIPE_system_input_pipe_188_inst_req_1 : boolean;
  signal RPIPE_system_input_pipe_188_inst_ack_1 : boolean;
  signal type_cast_192_inst_req_0 : boolean;
  signal type_cast_192_inst_ack_0 : boolean;
  signal type_cast_192_inst_req_1 : boolean;
  signal type_cast_192_inst_ack_1 : boolean;
  signal RPIPE_system_input_pipe_206_inst_req_0 : boolean;
  signal RPIPE_system_input_pipe_206_inst_ack_0 : boolean;
  signal RPIPE_system_input_pipe_206_inst_req_1 : boolean;
  signal RPIPE_system_input_pipe_206_inst_ack_1 : boolean;
  signal type_cast_210_inst_req_0 : boolean;
  signal type_cast_210_inst_ack_0 : boolean;
  signal type_cast_210_inst_req_1 : boolean;
  signal type_cast_210_inst_ack_1 : boolean;
  signal call_stmt_219_call_req_0 : boolean;
  signal call_stmt_219_call_ack_0 : boolean;
  signal call_stmt_219_call_req_1 : boolean;
  signal call_stmt_219_call_ack_1 : boolean;
  signal if_stmt_232_branch_req_0 : boolean;
  signal if_stmt_232_branch_ack_1 : boolean;
  signal if_stmt_232_branch_ack_0 : boolean;
  signal phi_stmt_76_req_0 : boolean;
  signal type_cast_82_inst_req_0 : boolean;
  signal type_cast_82_inst_ack_0 : boolean;
  signal type_cast_82_inst_req_1 : boolean;
  signal type_cast_82_inst_ack_1 : boolean;
  signal phi_stmt_76_req_1 : boolean;
  signal phi_stmt_76_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "fill_input_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  fill_input_CP_122_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "fill_input_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= fill_input_CP_122_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= fill_input_CP_122_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= fill_input_CP_122_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  fill_input_CP_122: Block -- control-path 
    signal fill_input_CP_122_elements: BooleanArray(43 downto 0);
    -- 
  begin -- 
    fill_input_CP_122_elements(0) <= fill_input_CP_122_start;
    fill_input_CP_122_symbol <= fill_input_CP_122_elements(36);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	38 
    -- CP-element group 0:  members (7) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_73/$entry
      -- CP-element group 0: 	 branch_block_stmt_73/branch_block_stmt_73__entry__
      -- CP-element group 0: 	 branch_block_stmt_73/bbx_xnph_forx_xbody
      -- CP-element group 0: 	 branch_block_stmt_73/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_73/bbx_xnph_forx_xbody_PhiReq/phi_stmt_76/$entry
      -- CP-element group 0: 	 branch_block_stmt_73/bbx_xnph_forx_xbody_PhiReq/phi_stmt_76/phi_stmt_76_sources/$entry
      -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	43 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_85_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_85_update_start_
      -- CP-element group 1: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_85_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_85_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_85_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_85_Update/cr
      -- 
    ra_151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_system_input_pipe_85_inst_ack_0, ack => fill_input_CP_122_elements(1)); -- 
    cr_155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(1), ack => RPIPE_system_input_pipe_85_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_85_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_85_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_85_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_89_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_89_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_89_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_98_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_98_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_98_Sample/rr
      -- 
    ca_156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_system_input_pipe_85_inst_ack_1, ack => fill_input_CP_122_elements(2)); -- 
    rr_164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(2), ack => type_cast_89_inst_req_0); -- 
    rr_178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(2), ack => RPIPE_system_input_pipe_98_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_89_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_89_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_89_Sample/ra
      -- 
    ra_165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_89_inst_ack_0, ack => fill_input_CP_122_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	43 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	33 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_89_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_89_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_89_Update/ca
      -- 
    ca_170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_89_inst_ack_1, ack => fill_input_CP_122_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_98_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_98_update_start_
      -- CP-element group 5: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_98_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_98_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_98_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_98_Update/cr
      -- 
    ra_179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_system_input_pipe_98_inst_ack_0, ack => fill_input_CP_122_elements(5)); -- 
    cr_183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(5), ack => RPIPE_system_input_pipe_98_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_98_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_98_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_98_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_102_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_102_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_102_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_116_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_116_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_116_Sample/rr
      -- 
    ca_184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_system_input_pipe_98_inst_ack_1, ack => fill_input_CP_122_elements(6)); -- 
    rr_192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(6), ack => type_cast_102_inst_req_0); -- 
    rr_206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(6), ack => RPIPE_system_input_pipe_116_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_102_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_102_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_102_Sample/ra
      -- 
    ra_193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_102_inst_ack_0, ack => fill_input_CP_122_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	43 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	33 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_102_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_102_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_102_Update/ca
      -- 
    ca_198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_102_inst_ack_1, ack => fill_input_CP_122_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_116_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_116_update_start_
      -- CP-element group 9: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_116_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_116_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_116_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_116_Update/cr
      -- 
    ra_207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_system_input_pipe_116_inst_ack_0, ack => fill_input_CP_122_elements(9)); -- 
    cr_211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(9), ack => RPIPE_system_input_pipe_116_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_116_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_116_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_116_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_120_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_120_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_120_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_134_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_134_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_134_Sample/rr
      -- 
    ca_212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_system_input_pipe_116_inst_ack_1, ack => fill_input_CP_122_elements(10)); -- 
    rr_220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(10), ack => type_cast_120_inst_req_0); -- 
    rr_234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(10), ack => RPIPE_system_input_pipe_134_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_120_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_120_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_120_Sample/ra
      -- 
    ra_221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_120_inst_ack_0, ack => fill_input_CP_122_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	43 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	33 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_120_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_120_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_120_Update/ca
      -- 
    ca_226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_120_inst_ack_1, ack => fill_input_CP_122_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_134_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_134_update_start_
      -- CP-element group 13: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_134_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_134_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_134_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_134_Update/cr
      -- 
    ra_235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_system_input_pipe_134_inst_ack_0, ack => fill_input_CP_122_elements(13)); -- 
    cr_239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(13), ack => RPIPE_system_input_pipe_134_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_138_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_152_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_152_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_134_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_134_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_134_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_138_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_138_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_152_Sample/rr
      -- 
    ca_240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_system_input_pipe_134_inst_ack_1, ack => fill_input_CP_122_elements(14)); -- 
    rr_248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(14), ack => type_cast_138_inst_req_0); -- 
    rr_262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(14), ack => RPIPE_system_input_pipe_152_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_138_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_138_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_138_Sample/$exit
      -- 
    ra_249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_138_inst_ack_0, ack => fill_input_CP_122_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	43 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	33 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_138_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_138_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_138_update_completed_
      -- 
    ca_254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_138_inst_ack_1, ack => fill_input_CP_122_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_152_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_152_update_start_
      -- CP-element group 17: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_152_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_152_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_152_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_152_Update/cr
      -- 
    ra_263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_system_input_pipe_152_inst_ack_0, ack => fill_input_CP_122_elements(17)); -- 
    cr_267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(17), ack => RPIPE_system_input_pipe_152_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_152_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_152_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_152_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_156_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_156_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_156_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_170_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_170_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_170_Sample/rr
      -- 
    ca_268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_system_input_pipe_152_inst_ack_1, ack => fill_input_CP_122_elements(18)); -- 
    rr_276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(18), ack => type_cast_156_inst_req_0); -- 
    rr_290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(18), ack => RPIPE_system_input_pipe_170_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_156_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_156_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_156_Sample/ra
      -- 
    ra_277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_156_inst_ack_0, ack => fill_input_CP_122_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	43 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	33 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_156_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_156_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_156_Update/ca
      -- 
    ca_282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_156_inst_ack_1, ack => fill_input_CP_122_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_170_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_170_update_start_
      -- CP-element group 21: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_170_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_170_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_170_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_170_Update/cr
      -- 
    ra_291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_system_input_pipe_170_inst_ack_0, ack => fill_input_CP_122_elements(21)); -- 
    cr_295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(21), ack => RPIPE_system_input_pipe_170_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_170_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_170_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_170_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_174_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_174_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_174_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_188_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_188_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_188_Sample/rr
      -- 
    ca_296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_system_input_pipe_170_inst_ack_1, ack => fill_input_CP_122_elements(22)); -- 
    rr_304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(22), ack => type_cast_174_inst_req_0); -- 
    rr_318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(22), ack => RPIPE_system_input_pipe_188_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_174_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_174_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_174_Sample/ra
      -- 
    ra_305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_174_inst_ack_0, ack => fill_input_CP_122_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	43 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	33 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_174_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_174_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_174_Update/ca
      -- 
    ca_310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_174_inst_ack_1, ack => fill_input_CP_122_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_188_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_188_update_start_
      -- CP-element group 25: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_188_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_188_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_188_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_188_Update/cr
      -- 
    ra_319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_system_input_pipe_188_inst_ack_0, ack => fill_input_CP_122_elements(25)); -- 
    cr_323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(25), ack => RPIPE_system_input_pipe_188_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_188_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_188_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_188_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_192_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_192_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_192_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_206_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_206_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_206_Sample/rr
      -- 
    ca_324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_system_input_pipe_188_inst_ack_1, ack => fill_input_CP_122_elements(26)); -- 
    rr_332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(26), ack => type_cast_192_inst_req_0); -- 
    rr_346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(26), ack => RPIPE_system_input_pipe_206_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_192_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_192_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_192_Sample/ra
      -- 
    ra_333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_192_inst_ack_0, ack => fill_input_CP_122_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	43 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	33 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_192_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_192_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_192_Update/ca
      -- 
    ca_338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_192_inst_ack_1, ack => fill_input_CP_122_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_206_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_206_update_start_
      -- CP-element group 29: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_206_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_206_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_206_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_206_Update/cr
      -- 
    ra_347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_system_input_pipe_206_inst_ack_0, ack => fill_input_CP_122_elements(29)); -- 
    cr_351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(29), ack => RPIPE_system_input_pipe_206_inst_req_1); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_206_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_206_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_206_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_210_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_210_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_210_Sample/rr
      -- 
    ca_352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_system_input_pipe_206_inst_ack_1, ack => fill_input_CP_122_elements(30)); -- 
    rr_360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(30), ack => type_cast_210_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_210_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_210_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_210_Sample/ra
      -- 
    ra_361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_210_inst_ack_0, ack => fill_input_CP_122_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	43 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_210_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_210_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_210_Update/ca
      -- 
    ca_366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_210_inst_ack_1, ack => fill_input_CP_122_elements(32)); -- 
    -- CP-element group 33:  join  transition  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	4 
    -- CP-element group 33: 	8 
    -- CP-element group 33: 	12 
    -- CP-element group 33: 	16 
    -- CP-element group 33: 	20 
    -- CP-element group 33: 	24 
    -- CP-element group 33: 	28 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/call_stmt_219_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/call_stmt_219_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/call_stmt_219_Sample/crr
      -- 
    crr_374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(33), ack => call_stmt_219_call_req_0); -- 
    fill_input_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 30) := "fill_input_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= fill_input_CP_122_elements(4) & fill_input_CP_122_elements(8) & fill_input_CP_122_elements(12) & fill_input_CP_122_elements(16) & fill_input_CP_122_elements(20) & fill_input_CP_122_elements(24) & fill_input_CP_122_elements(28) & fill_input_CP_122_elements(32);
      gj_fill_input_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_input_CP_122_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/call_stmt_219_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/call_stmt_219_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/call_stmt_219_Sample/cra
      -- 
    cra_375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_219_call_ack_0, ack => fill_input_CP_122_elements(34)); -- 
    -- CP-element group 35:  branch  transition  place  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	43 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (13) 
      -- CP-element group 35: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231__exit__
      -- CP-element group 35: 	 branch_block_stmt_73/if_stmt_232__entry__
      -- CP-element group 35: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/$exit
      -- CP-element group 35: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/call_stmt_219_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/call_stmt_219_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/call_stmt_219_Update/cca
      -- CP-element group 35: 	 branch_block_stmt_73/if_stmt_232_dead_link/$entry
      -- CP-element group 35: 	 branch_block_stmt_73/if_stmt_232_eval_test/$entry
      -- CP-element group 35: 	 branch_block_stmt_73/if_stmt_232_eval_test/$exit
      -- CP-element group 35: 	 branch_block_stmt_73/if_stmt_232_eval_test/branch_req
      -- CP-element group 35: 	 branch_block_stmt_73/R_exitcond1_233_place
      -- CP-element group 35: 	 branch_block_stmt_73/if_stmt_232_if_link/$entry
      -- CP-element group 35: 	 branch_block_stmt_73/if_stmt_232_else_link/$entry
      -- 
    cca_380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_219_call_ack_1, ack => fill_input_CP_122_elements(35)); -- 
    branch_req_388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(35), ack => if_stmt_232_branch_req_0); -- 
    -- CP-element group 36:  merge  transition  place  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (21) 
      -- CP-element group 36: 	 $exit
      -- CP-element group 36: 	 branch_block_stmt_73/$exit
      -- CP-element group 36: 	 branch_block_stmt_73/branch_block_stmt_73__exit__
      -- CP-element group 36: 	 branch_block_stmt_73/merge_stmt_238__exit__
      -- CP-element group 36: 	 branch_block_stmt_73/return__
      -- CP-element group 36: 	 branch_block_stmt_73/merge_stmt_240__exit__
      -- CP-element group 36: 	 branch_block_stmt_73/if_stmt_232_if_link/$exit
      -- CP-element group 36: 	 branch_block_stmt_73/if_stmt_232_if_link/if_choice_transition
      -- CP-element group 36: 	 branch_block_stmt_73/forx_xbody_forx_xend
      -- CP-element group 36: 	 branch_block_stmt_73/forx_xbody_forx_xend_PhiReq/$entry
      -- CP-element group 36: 	 branch_block_stmt_73/forx_xbody_forx_xend_PhiReq/$exit
      -- CP-element group 36: 	 branch_block_stmt_73/merge_stmt_238_PhiReqMerge
      -- CP-element group 36: 	 branch_block_stmt_73/merge_stmt_238_PhiAck/$entry
      -- CP-element group 36: 	 branch_block_stmt_73/merge_stmt_238_PhiAck/$exit
      -- CP-element group 36: 	 branch_block_stmt_73/merge_stmt_238_PhiAck/dummy
      -- CP-element group 36: 	 branch_block_stmt_73/return___PhiReq/$entry
      -- CP-element group 36: 	 branch_block_stmt_73/return___PhiReq/$exit
      -- CP-element group 36: 	 branch_block_stmt_73/merge_stmt_240_PhiReqMerge
      -- CP-element group 36: 	 branch_block_stmt_73/merge_stmt_240_PhiAck/$entry
      -- CP-element group 36: 	 branch_block_stmt_73/merge_stmt_240_PhiAck/$exit
      -- CP-element group 36: 	 branch_block_stmt_73/merge_stmt_240_PhiAck/dummy
      -- 
    if_choice_transition_393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_232_branch_ack_1, ack => fill_input_CP_122_elements(36)); -- 
    -- CP-element group 37:  fork  transition  place  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	40 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (12) 
      -- CP-element group 37: 	 branch_block_stmt_73/if_stmt_232_else_link/$exit
      -- CP-element group 37: 	 branch_block_stmt_73/if_stmt_232_else_link/else_choice_transition
      -- CP-element group 37: 	 branch_block_stmt_73/forx_xbody_forx_xbody
      -- CP-element group 37: 	 branch_block_stmt_73/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 37: 	 branch_block_stmt_73/forx_xbody_forx_xbody_PhiReq/phi_stmt_76/$entry
      -- CP-element group 37: 	 branch_block_stmt_73/forx_xbody_forx_xbody_PhiReq/phi_stmt_76/phi_stmt_76_sources/$entry
      -- CP-element group 37: 	 branch_block_stmt_73/forx_xbody_forx_xbody_PhiReq/phi_stmt_76/phi_stmt_76_sources/type_cast_82/$entry
      -- CP-element group 37: 	 branch_block_stmt_73/forx_xbody_forx_xbody_PhiReq/phi_stmt_76/phi_stmt_76_sources/type_cast_82/SplitProtocol/$entry
      -- CP-element group 37: 	 branch_block_stmt_73/forx_xbody_forx_xbody_PhiReq/phi_stmt_76/phi_stmt_76_sources/type_cast_82/SplitProtocol/Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_73/forx_xbody_forx_xbody_PhiReq/phi_stmt_76/phi_stmt_76_sources/type_cast_82/SplitProtocol/Sample/rr
      -- CP-element group 37: 	 branch_block_stmt_73/forx_xbody_forx_xbody_PhiReq/phi_stmt_76/phi_stmt_76_sources/type_cast_82/SplitProtocol/Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_73/forx_xbody_forx_xbody_PhiReq/phi_stmt_76/phi_stmt_76_sources/type_cast_82/SplitProtocol/Update/cr
      -- 
    else_choice_transition_397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_232_branch_ack_0, ack => fill_input_CP_122_elements(37)); -- 
    rr_429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(37), ack => type_cast_82_inst_req_0); -- 
    cr_434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(37), ack => type_cast_82_inst_req_1); -- 
    -- CP-element group 38:  transition  output  delay-element  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	0 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	42 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 branch_block_stmt_73/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 38: 	 branch_block_stmt_73/bbx_xnph_forx_xbody_PhiReq/phi_stmt_76/$exit
      -- CP-element group 38: 	 branch_block_stmt_73/bbx_xnph_forx_xbody_PhiReq/phi_stmt_76/phi_stmt_76_sources/$exit
      -- CP-element group 38: 	 branch_block_stmt_73/bbx_xnph_forx_xbody_PhiReq/phi_stmt_76/phi_stmt_76_sources/type_cast_80_konst_delay_trans
      -- CP-element group 38: 	 branch_block_stmt_73/bbx_xnph_forx_xbody_PhiReq/phi_stmt_76/phi_stmt_76_req
      -- 
    phi_stmt_76_req_410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_76_req_410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(38), ack => phi_stmt_76_req_0); -- 
    -- Element group fill_input_CP_122_elements(38) is a control-delay.
    cp_element_38_delay: control_delay_element  generic map(name => " 38_delay", delay_value => 1)  port map(req => fill_input_CP_122_elements(0), ack => fill_input_CP_122_elements(38), clk => clk, reset =>reset);
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_73/forx_xbody_forx_xbody_PhiReq/phi_stmt_76/phi_stmt_76_sources/type_cast_82/SplitProtocol/Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_73/forx_xbody_forx_xbody_PhiReq/phi_stmt_76/phi_stmt_76_sources/type_cast_82/SplitProtocol/Sample/ra
      -- 
    ra_430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_82_inst_ack_0, ack => fill_input_CP_122_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	37 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (2) 
      -- CP-element group 40: 	 branch_block_stmt_73/forx_xbody_forx_xbody_PhiReq/phi_stmt_76/phi_stmt_76_sources/type_cast_82/SplitProtocol/Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_73/forx_xbody_forx_xbody_PhiReq/phi_stmt_76/phi_stmt_76_sources/type_cast_82/SplitProtocol/Update/ca
      -- 
    ca_435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_82_inst_ack_1, ack => fill_input_CP_122_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_73/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 41: 	 branch_block_stmt_73/forx_xbody_forx_xbody_PhiReq/phi_stmt_76/$exit
      -- CP-element group 41: 	 branch_block_stmt_73/forx_xbody_forx_xbody_PhiReq/phi_stmt_76/phi_stmt_76_sources/$exit
      -- CP-element group 41: 	 branch_block_stmt_73/forx_xbody_forx_xbody_PhiReq/phi_stmt_76/phi_stmt_76_sources/type_cast_82/$exit
      -- CP-element group 41: 	 branch_block_stmt_73/forx_xbody_forx_xbody_PhiReq/phi_stmt_76/phi_stmt_76_sources/type_cast_82/SplitProtocol/$exit
      -- CP-element group 41: 	 branch_block_stmt_73/forx_xbody_forx_xbody_PhiReq/phi_stmt_76/phi_stmt_76_req
      -- 
    phi_stmt_76_req_436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_76_req_436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(41), ack => phi_stmt_76_req_1); -- 
    fill_input_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "fill_input_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_input_CP_122_elements(40) & fill_input_CP_122_elements(39);
      gj_fill_input_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_input_CP_122_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  merge  transition  place  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: 	38 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_73/merge_stmt_75_PhiReqMerge
      -- CP-element group 42: 	 branch_block_stmt_73/merge_stmt_75_PhiAck/$entry
      -- 
    fill_input_CP_122_elements(42) <= OrReduce(fill_input_CP_122_elements(41) & fill_input_CP_122_elements(38));
    -- CP-element group 43:  fork  transition  place  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	1 
    -- CP-element group 43: 	4 
    -- CP-element group 43: 	8 
    -- CP-element group 43: 	12 
    -- CP-element group 43: 	16 
    -- CP-element group 43: 	20 
    -- CP-element group 43: 	24 
    -- CP-element group 43: 	28 
    -- CP-element group 43: 	32 
    -- CP-element group 43: 	35 
    -- CP-element group 43:  members (35) 
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_138_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_138_Update/cr
      -- CP-element group 43: 	 branch_block_stmt_73/merge_stmt_75__exit__
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231__entry__
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/$entry
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_85_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_85_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/RPIPE_system_input_pipe_85_Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_89_update_start_
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_89_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_89_Update/cr
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_102_update_start_
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_102_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_102_Update/cr
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_120_update_start_
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_120_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_120_Update/cr
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_138_update_start_
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_156_update_start_
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_156_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_156_Update/cr
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_174_update_start_
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_174_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_174_Update/cr
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_192_update_start_
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_192_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_192_Update/cr
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_210_update_start_
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_210_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/type_cast_210_Update/cr
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/call_stmt_219_update_start_
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/call_stmt_219_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_73/assign_stmt_86_to_assign_stmt_231/call_stmt_219_Update/ccr
      -- CP-element group 43: 	 branch_block_stmt_73/merge_stmt_75_PhiAck/$exit
      -- CP-element group 43: 	 branch_block_stmt_73/merge_stmt_75_PhiAck/phi_stmt_76_ack
      -- 
    phi_stmt_76_ack_441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_76_ack_0, ack => fill_input_CP_122_elements(43)); -- 
    cr_253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(43), ack => type_cast_138_inst_req_1); -- 
    rr_150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(43), ack => RPIPE_system_input_pipe_85_inst_req_0); -- 
    cr_169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(43), ack => type_cast_89_inst_req_1); -- 
    cr_197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(43), ack => type_cast_102_inst_req_1); -- 
    cr_225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(43), ack => type_cast_120_inst_req_1); -- 
    cr_281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(43), ack => type_cast_156_inst_req_1); -- 
    cr_309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(43), ack => type_cast_174_inst_req_1); -- 
    cr_337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(43), ack => type_cast_192_inst_req_1); -- 
    cr_365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(43), ack => type_cast_210_inst_req_1); -- 
    ccr_379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_input_CP_122_elements(43), ack => call_stmt_219_call_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal add10_126 : std_logic_vector(63 downto 0);
    signal add16_144 : std_logic_vector(63 downto 0);
    signal add22_162 : std_logic_vector(63 downto 0);
    signal add28_180 : std_logic_vector(63 downto 0);
    signal add34_198 : std_logic_vector(63 downto 0);
    signal add40_216 : std_logic_vector(63 downto 0);
    signal add_108 : std_logic_vector(63 downto 0);
    signal call13_135 : std_logic_vector(7 downto 0);
    signal call19_153 : std_logic_vector(7 downto 0);
    signal call25_171 : std_logic_vector(7 downto 0);
    signal call2_99 : std_logic_vector(7 downto 0);
    signal call31_189 : std_logic_vector(7 downto 0);
    signal call37_207 : std_logic_vector(7 downto 0);
    signal call7_117 : std_logic_vector(7 downto 0);
    signal call_86 : std_logic_vector(7 downto 0);
    signal conv15_139 : std_logic_vector(63 downto 0);
    signal conv21_157 : std_logic_vector(63 downto 0);
    signal conv27_175 : std_logic_vector(63 downto 0);
    signal conv33_193 : std_logic_vector(63 downto 0);
    signal conv39_211 : std_logic_vector(63 downto 0);
    signal conv4_103 : std_logic_vector(63 downto 0);
    signal conv9_121 : std_logic_vector(63 downto 0);
    signal conv_90 : std_logic_vector(63 downto 0);
    signal exitcond1_231 : std_logic_vector(0 downto 0);
    signal iNsTr_1_76 : std_logic_vector(31 downto 0);
    signal inc_225 : std_logic_vector(31 downto 0);
    signal shl12_132 : std_logic_vector(63 downto 0);
    signal shl18_150 : std_logic_vector(63 downto 0);
    signal shl24_168 : std_logic_vector(63 downto 0);
    signal shl30_186 : std_logic_vector(63 downto 0);
    signal shl36_204 : std_logic_vector(63 downto 0);
    signal shl6_114 : std_logic_vector(63 downto 0);
    signal shl_96 : std_logic_vector(63 downto 0);
    signal type_cast_112_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_130_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_148_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_166_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_184_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_202_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_223_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_229_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_80_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_82_wire : std_logic_vector(31 downto 0);
    signal type_cast_94_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    type_cast_112_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_130_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_148_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_166_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_184_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_202_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_223_wire_constant <= "00000000000000000000000000000001";
    type_cast_229_wire_constant <= "00000000000000110001000000000000";
    type_cast_80_wire_constant <= "00000000000000000000000000000000";
    type_cast_94_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    phi_stmt_76: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_80_wire_constant & type_cast_82_wire;
      req <= phi_stmt_76_req_0 & phi_stmt_76_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_76",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_76_ack_0,
          idata => idata,
          odata => iNsTr_1_76,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_76
    type_cast_102_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_102_inst_req_0;
      type_cast_102_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_102_inst_req_1;
      type_cast_102_inst_ack_1<= rack(0);
      type_cast_102_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_102_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_99,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_120_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_120_inst_req_0;
      type_cast_120_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_120_inst_req_1;
      type_cast_120_inst_ack_1<= rack(0);
      type_cast_120_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_120_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call7_117,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9_121,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_138_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_138_inst_req_0;
      type_cast_138_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_138_inst_req_1;
      type_cast_138_inst_ack_1<= rack(0);
      type_cast_138_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_138_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call13_135,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv15_139,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_156_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_156_inst_req_0;
      type_cast_156_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_156_inst_req_1;
      type_cast_156_inst_ack_1<= rack(0);
      type_cast_156_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_156_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_153,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv21_157,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_174_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_174_inst_req_0;
      type_cast_174_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_174_inst_req_1;
      type_cast_174_inst_ack_1<= rack(0);
      type_cast_174_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_174_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call25_171,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv27_175,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_192_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_192_inst_req_0;
      type_cast_192_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_192_inst_req_1;
      type_cast_192_inst_ack_1<= rack(0);
      type_cast_192_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_192_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call31_189,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv33_193,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_210_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_210_inst_req_0;
      type_cast_210_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_210_inst_req_1;
      type_cast_210_inst_ack_1<= rack(0);
      type_cast_210_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_210_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_207,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_211,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_82_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_82_inst_req_0;
      type_cast_82_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_82_inst_req_1;
      type_cast_82_inst_ack_1<= rack(0);
      type_cast_82_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_82_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_225,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_82_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_89_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_89_inst_req_0;
      type_cast_89_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_89_inst_req_1;
      type_cast_89_inst_ack_1<= rack(0);
      type_cast_89_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_89_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_86,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_90,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    if_stmt_232_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_231;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_232_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_232_branch_req_0,
          ack0 => if_stmt_232_branch_ack_0,
          ack1 => if_stmt_232_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_224_inst
    process(iNsTr_1_76) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_1_76, type_cast_223_wire_constant, tmp_var);
      inc_225 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_230_inst
    process(inc_225) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_225, type_cast_229_wire_constant, tmp_var);
      exitcond1_231 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_107_inst
    process(shl_96, conv4_103) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_96, conv4_103, tmp_var);
      add_108 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_125_inst
    process(shl6_114, conv9_121) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl6_114, conv9_121, tmp_var);
      add10_126 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_143_inst
    process(shl12_132, conv15_139) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl12_132, conv15_139, tmp_var);
      add16_144 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_161_inst
    process(shl18_150, conv21_157) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_150, conv21_157, tmp_var);
      add22_162 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_179_inst
    process(shl24_168, conv27_175) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl24_168, conv27_175, tmp_var);
      add28_180 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_197_inst
    process(shl30_186, conv33_193) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl30_186, conv33_193, tmp_var);
      add34_198 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_215_inst
    process(shl36_204, conv39_211) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_204, conv39_211, tmp_var);
      add40_216 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_113_inst
    process(add_108) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add_108, type_cast_112_wire_constant, tmp_var);
      shl6_114 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_131_inst
    process(add10_126) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add10_126, type_cast_130_wire_constant, tmp_var);
      shl12_132 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_149_inst
    process(add16_144) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add16_144, type_cast_148_wire_constant, tmp_var);
      shl18_150 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_167_inst
    process(add22_162) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add22_162, type_cast_166_wire_constant, tmp_var);
      shl24_168 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_185_inst
    process(add28_180) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add28_180, type_cast_184_wire_constant, tmp_var);
      shl30_186 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_203_inst
    process(add34_198) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add34_198, type_cast_202_wire_constant, tmp_var);
      shl36_204 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_95_inst
    process(conv_90) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_90, type_cast_94_wire_constant, tmp_var);
      shl_96 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_system_input_pipe_85_inst RPIPE_system_input_pipe_98_inst RPIPE_system_input_pipe_116_inst RPIPE_system_input_pipe_134_inst RPIPE_system_input_pipe_152_inst RPIPE_system_input_pipe_170_inst RPIPE_system_input_pipe_188_inst RPIPE_system_input_pipe_206_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 7 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant outBUFs : IntegerArray(7 downto 0) := (7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      reqL_unguarded(7) <= RPIPE_system_input_pipe_85_inst_req_0;
      reqL_unguarded(6) <= RPIPE_system_input_pipe_98_inst_req_0;
      reqL_unguarded(5) <= RPIPE_system_input_pipe_116_inst_req_0;
      reqL_unguarded(4) <= RPIPE_system_input_pipe_134_inst_req_0;
      reqL_unguarded(3) <= RPIPE_system_input_pipe_152_inst_req_0;
      reqL_unguarded(2) <= RPIPE_system_input_pipe_170_inst_req_0;
      reqL_unguarded(1) <= RPIPE_system_input_pipe_188_inst_req_0;
      reqL_unguarded(0) <= RPIPE_system_input_pipe_206_inst_req_0;
      RPIPE_system_input_pipe_85_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_system_input_pipe_98_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_system_input_pipe_116_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_system_input_pipe_134_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_system_input_pipe_152_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_system_input_pipe_170_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_system_input_pipe_188_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_system_input_pipe_206_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= RPIPE_system_input_pipe_85_inst_req_1;
      reqR_unguarded(6) <= RPIPE_system_input_pipe_98_inst_req_1;
      reqR_unguarded(5) <= RPIPE_system_input_pipe_116_inst_req_1;
      reqR_unguarded(4) <= RPIPE_system_input_pipe_134_inst_req_1;
      reqR_unguarded(3) <= RPIPE_system_input_pipe_152_inst_req_1;
      reqR_unguarded(2) <= RPIPE_system_input_pipe_170_inst_req_1;
      reqR_unguarded(1) <= RPIPE_system_input_pipe_188_inst_req_1;
      reqR_unguarded(0) <= RPIPE_system_input_pipe_206_inst_req_1;
      RPIPE_system_input_pipe_85_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_system_input_pipe_98_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_system_input_pipe_116_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_system_input_pipe_134_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_system_input_pipe_152_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_system_input_pipe_170_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_system_input_pipe_188_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_system_input_pipe_206_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      call_86 <= data_out(63 downto 56);
      call2_99 <= data_out(55 downto 48);
      call7_117 <= data_out(47 downto 40);
      call13_135 <= data_out(39 downto 32);
      call19_153 <= data_out(31 downto 24);
      call25_171 <= data_out(23 downto 16);
      call31_189 <= data_out(15 downto 8);
      call37_207 <= data_out(7 downto 0);
      system_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "system_input_pipe_read_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      system_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "system_input_pipe_read_0", data_width => 8,  num_reqs => 8,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => system_input_pipe_pipe_read_req(0),
          oack => system_input_pipe_pipe_read_ack(0),
          odata => system_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared call operator group (0) : call_stmt_219_call 
    writeModule1_call_group_0: Block -- 
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_219_call_req_0;
      call_stmt_219_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_219_call_req_1;
      call_stmt_219_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writeModule1_call_group_0_gI: SplitGuardInterface generic map(name => "writeModule1_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= iNsTr_1_76 & add40_216;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 96,
        owidth => 96,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writeModule1_call_reqs(0),
          ackR => writeModule1_call_acks(0),
          dataR => writeModule1_call_data(95 downto 0),
          tagR => writeModule1_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => writeModule1_return_acks(0), -- cross-over
          ackL => writeModule1_return_reqs(0), -- cross-over
          tagL => writeModule1_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end fill_input_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity maxPool4 is -- 
  generic (tag_length : integer); 
  port ( -- 
    addr : in  std_logic_vector(31 downto 0);
    addr1 : in  std_logic_vector(31 downto 0);
    addr2 : in  std_logic_vector(31 downto 0);
    addr3 : in  std_logic_vector(31 downto 0);
    addr4 : in  std_logic_vector(31 downto 0);
    index1 : in  std_logic_vector(7 downto 0);
    index2 : in  std_logic_vector(7 downto 0);
    output : out  std_logic_vector(7 downto 0);
    readModule_maxPool_call_reqs : out  std_logic_vector(0 downto 0);
    readModule_maxPool_call_acks : in   std_logic_vector(0 downto 0);
    readModule_maxPool_call_data : out  std_logic_vector(39 downto 0);
    readModule_maxPool_call_tag  :  out  std_logic_vector(2 downto 0);
    readModule_maxPool_return_reqs : out  std_logic_vector(0 downto 0);
    readModule_maxPool_return_acks : in   std_logic_vector(0 downto 0);
    readModule_maxPool_return_data : in   std_logic_vector(63 downto 0);
    readModule_maxPool_return_tag :  in   std_logic_vector(2 downto 0);
    writeModule_maxPool_call_reqs : out  std_logic_vector(0 downto 0);
    writeModule_maxPool_call_acks : in   std_logic_vector(0 downto 0);
    writeModule_maxPool_call_data : out  std_logic_vector(103 downto 0);
    writeModule_maxPool_call_tag  :  out  std_logic_vector(0 downto 0);
    writeModule_maxPool_return_reqs : out  std_logic_vector(0 downto 0);
    writeModule_maxPool_return_acks : in   std_logic_vector(0 downto 0);
    writeModule_maxPool_return_data : in   std_logic_vector(0 downto 0);
    writeModule_maxPool_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity maxPool4;
architecture maxPool4_arch of maxPool4 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 176)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal addr_buffer :  std_logic_vector(31 downto 0);
  signal addr_update_enable: Boolean;
  signal addr1_buffer :  std_logic_vector(31 downto 0);
  signal addr1_update_enable: Boolean;
  signal addr2_buffer :  std_logic_vector(31 downto 0);
  signal addr2_update_enable: Boolean;
  signal addr3_buffer :  std_logic_vector(31 downto 0);
  signal addr3_update_enable: Boolean;
  signal addr4_buffer :  std_logic_vector(31 downto 0);
  signal addr4_update_enable: Boolean;
  signal index1_buffer :  std_logic_vector(7 downto 0);
  signal index1_update_enable: Boolean;
  signal index2_buffer :  std_logic_vector(7 downto 0);
  signal index2_update_enable: Boolean;
  -- output port buffer signals
  signal output_buffer :  std_logic_vector(7 downto 0);
  signal output_update_enable: Boolean;
  signal maxPool4_CP_563_start: Boolean;
  signal maxPool4_CP_563_symbol: Boolean;
  -- volatile/operator module components. 
  component readModule_maxPool is -- 
    generic (tag_length : integer); 
    port ( -- 
      index : in  std_logic_vector(7 downto 0);
      address : in  std_logic_vector(31 downto 0);
      data : out  std_logic_vector(63 downto 0);
      memoryModule_call_reqs : out  std_logic_vector(0 downto 0);
      memoryModule_call_acks : in   std_logic_vector(0 downto 0);
      memoryModule_call_data : out  std_logic_vector(96 downto 0);
      memoryModule_call_tag  :  out  std_logic_vector(0 downto 0);
      memoryModule_return_reqs : out  std_logic_vector(0 downto 0);
      memoryModule_return_acks : in   std_logic_vector(0 downto 0);
      memoryModule_return_data : in   std_logic_vector(63 downto 0);
      memoryModule_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component writeModule_maxPool is -- 
    generic (tag_length : integer); 
    port ( -- 
      index : in  std_logic_vector(7 downto 0);
      address : in  std_logic_vector(31 downto 0);
      data : in  std_logic_vector(63 downto 0);
      done : out  std_logic_vector(0 downto 0);
      memoryModule_call_reqs : out  std_logic_vector(0 downto 0);
      memoryModule_call_acks : in   std_logic_vector(0 downto 0);
      memoryModule_call_data : out  std_logic_vector(96 downto 0);
      memoryModule_call_tag  :  out  std_logic_vector(0 downto 0);
      memoryModule_return_reqs : out  std_logic_vector(0 downto 0);
      memoryModule_return_acks : in   std_logic_vector(0 downto 0);
      memoryModule_return_data : in   std_logic_vector(63 downto 0);
      memoryModule_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal slice_344_inst_ack_1 : boolean;
  signal slice_332_inst_req_1 : boolean;
  signal slice_344_inst_req_0 : boolean;
  signal slice_344_inst_ack_0 : boolean;
  signal slice_344_inst_req_1 : boolean;
  signal slice_308_inst_ack_1 : boolean;
  signal slice_308_inst_req_1 : boolean;
  signal slice_320_inst_req_1 : boolean;
  signal call_stmt_305_call_ack_1 : boolean;
  signal slice_308_inst_ack_0 : boolean;
  signal slice_336_inst_ack_0 : boolean;
  signal slice_308_inst_req_0 : boolean;
  signal slice_320_inst_ack_0 : boolean;
  signal call_stmt_301_call_ack_1 : boolean;
  signal slice_332_inst_ack_0 : boolean;
  signal slice_332_inst_req_0 : boolean;
  signal slice_316_inst_ack_1 : boolean;
  signal slice_336_inst_req_0 : boolean;
  signal call_stmt_305_call_req_1 : boolean;
  signal slice_316_inst_ack_0 : boolean;
  signal slice_332_inst_ack_1 : boolean;
  signal slice_316_inst_req_0 : boolean;
  signal slice_312_inst_req_1 : boolean;
  signal slice_316_inst_req_1 : boolean;
  signal call_stmt_301_call_req_1 : boolean;
  signal call_stmt_305_call_ack_0 : boolean;
  signal slice_320_inst_req_0 : boolean;
  signal call_stmt_293_call_ack_1 : boolean;
  signal call_stmt_305_call_req_0 : boolean;
  signal call_stmt_293_call_req_1 : boolean;
  signal call_stmt_293_call_ack_0 : boolean;
  signal slice_348_inst_req_0 : boolean;
  signal slice_348_inst_ack_0 : boolean;
  signal slice_312_inst_ack_1 : boolean;
  signal slice_356_inst_req_1 : boolean;
  signal slice_356_inst_ack_1 : boolean;
  signal call_stmt_301_call_ack_0 : boolean;
  signal call_stmt_293_call_req_0 : boolean;
  signal slice_312_inst_ack_0 : boolean;
  signal call_stmt_301_call_req_0 : boolean;
  signal slice_312_inst_req_0 : boolean;
  signal call_stmt_297_call_ack_1 : boolean;
  signal call_stmt_297_call_req_1 : boolean;
  signal call_stmt_297_call_ack_0 : boolean;
  signal call_stmt_297_call_req_0 : boolean;
  signal slice_340_inst_req_0 : boolean;
  signal slice_336_inst_req_1 : boolean;
  signal slice_320_inst_ack_1 : boolean;
  signal slice_328_inst_ack_1 : boolean;
  signal slice_328_inst_req_1 : boolean;
  signal slice_328_inst_ack_0 : boolean;
  signal slice_328_inst_req_0 : boolean;
  signal slice_324_inst_ack_1 : boolean;
  signal slice_324_inst_req_1 : boolean;
  signal slice_336_inst_ack_1 : boolean;
  signal slice_340_inst_ack_1 : boolean;
  signal slice_340_inst_req_1 : boolean;
  signal slice_340_inst_ack_0 : boolean;
  signal slice_348_inst_req_1 : boolean;
  signal slice_348_inst_ack_1 : boolean;
  signal slice_352_inst_req_0 : boolean;
  signal slice_356_inst_req_0 : boolean;
  signal slice_324_inst_ack_0 : boolean;
  signal slice_324_inst_req_0 : boolean;
  signal slice_356_inst_ack_0 : boolean;
  signal slice_352_inst_req_1 : boolean;
  signal slice_352_inst_ack_1 : boolean;
  signal slice_352_inst_ack_0 : boolean;
  signal slice_360_inst_req_0 : boolean;
  signal slice_360_inst_ack_0 : boolean;
  signal slice_360_inst_req_1 : boolean;
  signal slice_360_inst_ack_1 : boolean;
  signal slice_364_inst_req_0 : boolean;
  signal slice_364_inst_ack_0 : boolean;
  signal slice_364_inst_req_1 : boolean;
  signal slice_364_inst_ack_1 : boolean;
  signal slice_368_inst_req_0 : boolean;
  signal slice_368_inst_ack_0 : boolean;
  signal slice_368_inst_req_1 : boolean;
  signal slice_368_inst_ack_1 : boolean;
  signal slice_372_inst_req_0 : boolean;
  signal slice_372_inst_ack_0 : boolean;
  signal slice_372_inst_req_1 : boolean;
  signal slice_372_inst_ack_1 : boolean;
  signal slice_376_inst_req_0 : boolean;
  signal slice_376_inst_ack_0 : boolean;
  signal slice_376_inst_req_1 : boolean;
  signal slice_376_inst_ack_1 : boolean;
  signal slice_380_inst_req_0 : boolean;
  signal slice_380_inst_ack_0 : boolean;
  signal slice_380_inst_req_1 : boolean;
  signal slice_380_inst_ack_1 : boolean;
  signal slice_384_inst_req_0 : boolean;
  signal slice_384_inst_ack_0 : boolean;
  signal slice_384_inst_req_1 : boolean;
  signal slice_384_inst_ack_1 : boolean;
  signal slice_388_inst_req_0 : boolean;
  signal slice_388_inst_ack_0 : boolean;
  signal slice_388_inst_req_1 : boolean;
  signal slice_388_inst_ack_1 : boolean;
  signal slice_392_inst_req_0 : boolean;
  signal slice_392_inst_ack_0 : boolean;
  signal slice_392_inst_req_1 : boolean;
  signal slice_392_inst_ack_1 : boolean;
  signal slice_396_inst_req_0 : boolean;
  signal slice_396_inst_ack_0 : boolean;
  signal slice_396_inst_req_1 : boolean;
  signal slice_396_inst_ack_1 : boolean;
  signal slice_400_inst_req_0 : boolean;
  signal slice_400_inst_ack_0 : boolean;
  signal slice_400_inst_req_1 : boolean;
  signal slice_400_inst_ack_1 : boolean;
  signal slice_404_inst_req_0 : boolean;
  signal slice_404_inst_ack_0 : boolean;
  signal slice_404_inst_req_1 : boolean;
  signal slice_404_inst_ack_1 : boolean;
  signal slice_408_inst_req_0 : boolean;
  signal slice_408_inst_ack_0 : boolean;
  signal slice_408_inst_req_1 : boolean;
  signal slice_408_inst_ack_1 : boolean;
  signal slice_412_inst_req_0 : boolean;
  signal slice_412_inst_ack_0 : boolean;
  signal slice_412_inst_req_1 : boolean;
  signal slice_412_inst_ack_1 : boolean;
  signal slice_416_inst_req_0 : boolean;
  signal slice_416_inst_ack_0 : boolean;
  signal slice_416_inst_req_1 : boolean;
  signal slice_416_inst_ack_1 : boolean;
  signal slice_420_inst_req_0 : boolean;
  signal slice_420_inst_ack_0 : boolean;
  signal slice_420_inst_req_1 : boolean;
  signal slice_420_inst_ack_1 : boolean;
  signal slice_424_inst_req_0 : boolean;
  signal slice_424_inst_ack_0 : boolean;
  signal slice_424_inst_req_1 : boolean;
  signal slice_424_inst_ack_1 : boolean;
  signal slice_428_inst_req_0 : boolean;
  signal slice_428_inst_ack_0 : boolean;
  signal slice_428_inst_req_1 : boolean;
  signal slice_428_inst_ack_1 : boolean;
  signal slice_432_inst_req_0 : boolean;
  signal slice_432_inst_ack_0 : boolean;
  signal slice_432_inst_req_1 : boolean;
  signal slice_432_inst_ack_1 : boolean;
  signal W_index2_755_delayed_7_0_755_inst_req_0 : boolean;
  signal W_index2_755_delayed_7_0_755_inst_ack_0 : boolean;
  signal W_index2_755_delayed_7_0_755_inst_req_1 : boolean;
  signal W_index2_755_delayed_7_0_755_inst_ack_1 : boolean;
  signal W_addr_756_delayed_7_0_758_inst_req_0 : boolean;
  signal W_addr_756_delayed_7_0_758_inst_ack_0 : boolean;
  signal W_addr_756_delayed_7_0_758_inst_req_1 : boolean;
  signal W_addr_756_delayed_7_0_758_inst_ack_1 : boolean;
  signal call_stmt_788_call_req_0 : boolean;
  signal call_stmt_788_call_ack_0 : boolean;
  signal call_stmt_788_call_req_1 : boolean;
  signal call_stmt_788_call_ack_1 : boolean;
  signal type_cast_791_inst_req_0 : boolean;
  signal type_cast_791_inst_ack_0 : boolean;
  signal type_cast_791_inst_req_1 : boolean;
  signal type_cast_791_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "maxPool4_input_buffer", -- 
      buffer_size => 2,
      bypass_flag => false,
      data_width => tag_length + 176) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= addr;
  addr_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= addr1;
  addr1_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(95 downto 64) <= addr2;
  addr2_buffer <= in_buffer_data_out(95 downto 64);
  in_buffer_data_in(127 downto 96) <= addr3;
  addr3_buffer <= in_buffer_data_out(127 downto 96);
  in_buffer_data_in(159 downto 128) <= addr4;
  addr4_buffer <= in_buffer_data_out(159 downto 128);
  in_buffer_data_in(167 downto 160) <= index1;
  index1_buffer <= in_buffer_data_out(167 downto 160);
  in_buffer_data_in(175 downto 168) <= index2;
  index2_buffer <= in_buffer_data_out(175 downto 168);
  in_buffer_data_in(tag_length + 175 downto 176) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 175 downto 176);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 8) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 1,8 => 15);
    constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1,8 => 15);
    constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 9); -- 
  begin -- 
    preds <= addr_update_enable & addr1_update_enable & addr2_update_enable & addr3_update_enable & addr4_update_enable & index1_update_enable & index2_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  maxPool4_CP_563_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "maxPool4_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= output_buffer;
  output <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 15);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool4_CP_563_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  output_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 25) := "output_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_output_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => output_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 15,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= maxPool4_CP_563_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool4_CP_563_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  maxPool4_CP_563: Block -- control-path 
    signal maxPool4_CP_563_elements: BooleanArray(179 downto 0);
    -- 
  begin -- 
    maxPool4_CP_563_elements(0) <= maxPool4_CP_563_start;
    maxPool4_CP_563_symbol <= maxPool4_CP_563_elements(179);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	10 
    -- CP-element group 1: 	18 
    -- CP-element group 1: 	22 
    -- CP-element group 1: 	14 
    -- CP-element group 1: 	154 
    -- CP-element group 1: 	158 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 call_stmt_293_to_assign_stmt_792/$entry
      -- 
    maxPool4_CP_563_elements(1) <= maxPool4_CP_563_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	160 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	171 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 call_stmt_293_to_assign_stmt_792/addr_update_enable
      -- CP-element group 2: 	 call_stmt_293_to_assign_stmt_792/addr_update_enable_out
      -- 
    maxPool4_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_563_elements(160);
      gj_maxPool4_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	12 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	172 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 call_stmt_293_to_assign_stmt_792/addr1_update_enable_out
      -- CP-element group 3: 	 call_stmt_293_to_assign_stmt_792/addr1_update_enable
      -- 
    maxPool4_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_563_elements(12);
      gj_maxPool4_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	16 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	173 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 call_stmt_293_to_assign_stmt_792/addr2_update_enable_out
      -- CP-element group 4: 	 call_stmt_293_to_assign_stmt_792/addr2_update_enable
      -- 
    maxPool4_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_563_elements(16);
      gj_maxPool4_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	20 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	174 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 call_stmt_293_to_assign_stmt_792/addr3_update_enable_out
      -- CP-element group 5: 	 call_stmt_293_to_assign_stmt_792/addr3_update_enable
      -- 
    maxPool4_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_563_elements(20);
      gj_maxPool4_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	24 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	175 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 call_stmt_293_to_assign_stmt_792/addr4_update_enable_out
      -- CP-element group 6: 	 call_stmt_293_to_assign_stmt_792/addr4_update_enable
      -- 
    maxPool4_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_563_elements(24);
      gj_maxPool4_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  join  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: marked-predecessors 
    -- CP-element group 7: 	12 
    -- CP-element group 7: 	16 
    -- CP-element group 7: 	20 
    -- CP-element group 7: 	24 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	176 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 call_stmt_293_to_assign_stmt_792/index1_update_enable_out
      -- CP-element group 7: 	 call_stmt_293_to_assign_stmt_792/index1_update_enable
      -- 
    maxPool4_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(12) & maxPool4_CP_563_elements(16) & maxPool4_CP_563_elements(20) & maxPool4_CP_563_elements(24);
      gj_maxPool4_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  join  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	156 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	177 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 call_stmt_293_to_assign_stmt_792/index2_update_enable_out
      -- CP-element group 8: 	 call_stmt_293_to_assign_stmt_792/index2_update_enable
      -- 
    maxPool4_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_563_elements(156);
      gj_maxPool4_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	178 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	167 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 call_stmt_293_to_assign_stmt_792/output_update_enable_in
      -- CP-element group 9: 	 call_stmt_293_to_assign_stmt_792/output_update_enable
      -- 
    maxPool4_CP_563_elements(9) <= maxPool4_CP_563_elements(178);
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	1 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_293_to_assign_stmt_792/call_stmt_293_Sample/crr
      -- CP-element group 10: 	 call_stmt_293_to_assign_stmt_792/call_stmt_293_Sample/$entry
      -- CP-element group 10: 	 call_stmt_293_to_assign_stmt_792/call_stmt_293_sample_start_
      -- 
    crr_592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(10), ack => call_stmt_293_call_req_0); -- 
    maxPool4_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(1) & maxPool4_CP_563_elements(12);
      gj_maxPool4_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	40 
    -- CP-element group 11: 	44 
    -- CP-element group 11: 	48 
    -- CP-element group 11: 	52 
    -- CP-element group 11: 	56 
    -- CP-element group 11: 	13 
    -- CP-element group 11: 	28 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	32 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_293_to_assign_stmt_792/call_stmt_293_Update/ccr
      -- CP-element group 11: 	 call_stmt_293_to_assign_stmt_792/call_stmt_293_Update/$entry
      -- CP-element group 11: 	 call_stmt_293_to_assign_stmt_792/call_stmt_293_update_start_
      -- 
    ccr_597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(11), ack => call_stmt_293_call_req_1); -- 
    maxPool4_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(40) & maxPool4_CP_563_elements(44) & maxPool4_CP_563_elements(48) & maxPool4_CP_563_elements(52) & maxPool4_CP_563_elements(56) & maxPool4_CP_563_elements(13) & maxPool4_CP_563_elements(28) & maxPool4_CP_563_elements(36) & maxPool4_CP_563_elements(32);
      gj_maxPool4_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	7 
    -- CP-element group 12: 	3 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_293_to_assign_stmt_792/call_stmt_293_Sample/cra
      -- CP-element group 12: 	 call_stmt_293_to_assign_stmt_792/call_stmt_293_Sample/$exit
      -- CP-element group 12: 	 call_stmt_293_to_assign_stmt_792/call_stmt_293_sample_completed_
      -- 
    cra_593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_293_call_ack_0, ack => maxPool4_CP_563_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	42 
    -- CP-element group 13: 	46 
    -- CP-element group 13: 	50 
    -- CP-element group 13: 	54 
    -- CP-element group 13: 	26 
    -- CP-element group 13: 	34 
    -- CP-element group 13: 	30 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	11 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_293_to_assign_stmt_792/call_stmt_293_Update/cca
      -- CP-element group 13: 	 call_stmt_293_to_assign_stmt_792/call_stmt_293_Update/$exit
      -- CP-element group 13: 	 call_stmt_293_to_assign_stmt_792/call_stmt_293_update_completed_
      -- 
    cca_598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_293_call_ack_1, ack => maxPool4_CP_563_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	1 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 call_stmt_293_to_assign_stmt_792/call_stmt_297_Sample/$entry
      -- CP-element group 14: 	 call_stmt_293_to_assign_stmt_792/call_stmt_297_sample_start_
      -- CP-element group 14: 	 call_stmt_293_to_assign_stmt_792/call_stmt_297_Sample/crr
      -- 
    crr_606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(14), ack => call_stmt_297_call_req_0); -- 
    maxPool4_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(1) & maxPool4_CP_563_elements(16);
      gj_maxPool4_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	60 
    -- CP-element group 15: 	64 
    -- CP-element group 15: 	68 
    -- CP-element group 15: 	72 
    -- CP-element group 15: 	76 
    -- CP-element group 15: 	80 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	84 
    -- CP-element group 15: 	88 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 call_stmt_293_to_assign_stmt_792/call_stmt_297_update_start_
      -- CP-element group 15: 	 call_stmt_293_to_assign_stmt_792/call_stmt_297_Update/ccr
      -- CP-element group 15: 	 call_stmt_293_to_assign_stmt_792/call_stmt_297_Update/$entry
      -- 
    ccr_611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(15), ack => call_stmt_297_call_req_1); -- 
    maxPool4_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(60) & maxPool4_CP_563_elements(64) & maxPool4_CP_563_elements(68) & maxPool4_CP_563_elements(72) & maxPool4_CP_563_elements(76) & maxPool4_CP_563_elements(80) & maxPool4_CP_563_elements(17) & maxPool4_CP_563_elements(84) & maxPool4_CP_563_elements(88);
      gj_maxPool4_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	4 
    -- CP-element group 16: 	7 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 call_stmt_293_to_assign_stmt_792/call_stmt_297_sample_completed_
      -- CP-element group 16: 	 call_stmt_293_to_assign_stmt_792/call_stmt_297_Sample/cra
      -- CP-element group 16: 	 call_stmt_293_to_assign_stmt_792/call_stmt_297_Sample/$exit
      -- 
    cra_607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_297_call_ack_0, ack => maxPool4_CP_563_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	58 
    -- CP-element group 17: 	62 
    -- CP-element group 17: 	66 
    -- CP-element group 17: 	70 
    -- CP-element group 17: 	74 
    -- CP-element group 17: 	78 
    -- CP-element group 17: 	82 
    -- CP-element group 17: 	86 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	15 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 call_stmt_293_to_assign_stmt_792/call_stmt_297_update_completed_
      -- CP-element group 17: 	 call_stmt_293_to_assign_stmt_792/call_stmt_297_Update/cca
      -- CP-element group 17: 	 call_stmt_293_to_assign_stmt_792/call_stmt_297_Update/$exit
      -- 
    cca_612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_297_call_ack_1, ack => maxPool4_CP_563_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	1 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 call_stmt_293_to_assign_stmt_792/call_stmt_301_sample_start_
      -- CP-element group 18: 	 call_stmt_293_to_assign_stmt_792/call_stmt_301_Sample/crr
      -- CP-element group 18: 	 call_stmt_293_to_assign_stmt_792/call_stmt_301_Sample/$entry
      -- 
    crr_620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(18), ack => call_stmt_301_call_req_0); -- 
    maxPool4_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(1) & maxPool4_CP_563_elements(20);
      gj_maxPool4_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	21 
    -- CP-element group 19: 	92 
    -- CP-element group 19: 	96 
    -- CP-element group 19: 	100 
    -- CP-element group 19: 	104 
    -- CP-element group 19: 	108 
    -- CP-element group 19: 	112 
    -- CP-element group 19: 	116 
    -- CP-element group 19: 	120 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 call_stmt_293_to_assign_stmt_792/call_stmt_301_update_start_
      -- CP-element group 19: 	 call_stmt_293_to_assign_stmt_792/call_stmt_301_Update/ccr
      -- CP-element group 19: 	 call_stmt_293_to_assign_stmt_792/call_stmt_301_Update/$entry
      -- 
    ccr_625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(19), ack => call_stmt_301_call_req_1); -- 
    maxPool4_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(21) & maxPool4_CP_563_elements(92) & maxPool4_CP_563_elements(96) & maxPool4_CP_563_elements(100) & maxPool4_CP_563_elements(104) & maxPool4_CP_563_elements(108) & maxPool4_CP_563_elements(112) & maxPool4_CP_563_elements(116) & maxPool4_CP_563_elements(120);
      gj_maxPool4_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	7 
    -- CP-element group 20: 	18 
    -- CP-element group 20: 	5 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 call_stmt_293_to_assign_stmt_792/call_stmt_301_sample_completed_
      -- CP-element group 20: 	 call_stmt_293_to_assign_stmt_792/call_stmt_301_Sample/cra
      -- CP-element group 20: 	 call_stmt_293_to_assign_stmt_792/call_stmt_301_Sample/$exit
      -- 
    cra_621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_301_call_ack_0, ack => maxPool4_CP_563_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	90 
    -- CP-element group 21: 	94 
    -- CP-element group 21: 	98 
    -- CP-element group 21: 	102 
    -- CP-element group 21: 	106 
    -- CP-element group 21: 	110 
    -- CP-element group 21: 	114 
    -- CP-element group 21: 	118 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	19 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 call_stmt_293_to_assign_stmt_792/call_stmt_301_update_completed_
      -- CP-element group 21: 	 call_stmt_293_to_assign_stmt_792/call_stmt_301_Update/cca
      -- CP-element group 21: 	 call_stmt_293_to_assign_stmt_792/call_stmt_301_Update/$exit
      -- 
    cca_626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_301_call_ack_1, ack => maxPool4_CP_563_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	1 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 call_stmt_293_to_assign_stmt_792/call_stmt_305_sample_start_
      -- CP-element group 22: 	 call_stmt_293_to_assign_stmt_792/call_stmt_305_Sample/crr
      -- CP-element group 22: 	 call_stmt_293_to_assign_stmt_792/call_stmt_305_Sample/$entry
      -- 
    crr_634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(22), ack => call_stmt_305_call_req_0); -- 
    maxPool4_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(1) & maxPool4_CP_563_elements(24);
      gj_maxPool4_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: 	124 
    -- CP-element group 23: 	128 
    -- CP-element group 23: 	132 
    -- CP-element group 23: 	136 
    -- CP-element group 23: 	140 
    -- CP-element group 23: 	144 
    -- CP-element group 23: 	148 
    -- CP-element group 23: 	152 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 call_stmt_293_to_assign_stmt_792/call_stmt_305_Update/ccr
      -- CP-element group 23: 	 call_stmt_293_to_assign_stmt_792/call_stmt_305_Update/$entry
      -- CP-element group 23: 	 call_stmt_293_to_assign_stmt_792/call_stmt_305_update_start_
      -- 
    ccr_639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(23), ack => call_stmt_305_call_req_1); -- 
    maxPool4_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(25) & maxPool4_CP_563_elements(124) & maxPool4_CP_563_elements(128) & maxPool4_CP_563_elements(132) & maxPool4_CP_563_elements(136) & maxPool4_CP_563_elements(140) & maxPool4_CP_563_elements(144) & maxPool4_CP_563_elements(148) & maxPool4_CP_563_elements(152);
      gj_maxPool4_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	7 
    -- CP-element group 24: 	6 
    -- CP-element group 24: 	22 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 call_stmt_293_to_assign_stmt_792/call_stmt_305_Sample/cra
      -- CP-element group 24: 	 call_stmt_293_to_assign_stmt_792/call_stmt_305_Sample/$exit
      -- CP-element group 24: 	 call_stmt_293_to_assign_stmt_792/call_stmt_305_sample_completed_
      -- 
    cra_635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_305_call_ack_0, ack => maxPool4_CP_563_elements(24)); -- 
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	122 
    -- CP-element group 25: 	126 
    -- CP-element group 25: 	130 
    -- CP-element group 25: 	134 
    -- CP-element group 25: 	138 
    -- CP-element group 25: 	142 
    -- CP-element group 25: 	146 
    -- CP-element group 25: 	150 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	23 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 call_stmt_293_to_assign_stmt_792/call_stmt_305_Update/cca
      -- CP-element group 25: 	 call_stmt_293_to_assign_stmt_792/call_stmt_305_Update/$exit
      -- CP-element group 25: 	 call_stmt_293_to_assign_stmt_792/call_stmt_305_update_completed_
      -- 
    cca_640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_305_call_ack_1, ack => maxPool4_CP_563_elements(25)); -- 
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	13 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 call_stmt_293_to_assign_stmt_792/slice_308_Sample/rr
      -- CP-element group 26: 	 call_stmt_293_to_assign_stmt_792/slice_308_Sample/$entry
      -- CP-element group 26: 	 call_stmt_293_to_assign_stmt_792/slice_308_sample_start_
      -- 
    rr_648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(26), ack => slice_308_inst_req_0); -- 
    maxPool4_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(13) & maxPool4_CP_563_elements(28);
      gj_maxPool4_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: 	164 
    -- CP-element group 27: 	168 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 call_stmt_293_to_assign_stmt_792/slice_308_Update/cr
      -- CP-element group 27: 	 call_stmt_293_to_assign_stmt_792/slice_308_Update/$entry
      -- CP-element group 27: 	 call_stmt_293_to_assign_stmt_792/slice_308_update_start_
      -- 
    cr_653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(27), ack => slice_308_inst_req_1); -- 
    maxPool4_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(29) & maxPool4_CP_563_elements(164) & maxPool4_CP_563_elements(168);
      gj_maxPool4_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	11 
    -- CP-element group 28: 	26 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 call_stmt_293_to_assign_stmt_792/slice_308_Sample/ra
      -- CP-element group 28: 	 call_stmt_293_to_assign_stmt_792/slice_308_Sample/$exit
      -- CP-element group 28: 	 call_stmt_293_to_assign_stmt_792/slice_308_sample_completed_
      -- 
    ra_649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_308_inst_ack_0, ack => maxPool4_CP_563_elements(28)); -- 
    -- CP-element group 29:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	162 
    -- CP-element group 29: 	166 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 call_stmt_293_to_assign_stmt_792/slice_308_Update/ca
      -- CP-element group 29: 	 call_stmt_293_to_assign_stmt_792/slice_308_Update/$exit
      -- CP-element group 29: 	 call_stmt_293_to_assign_stmt_792/slice_308_update_completed_
      -- 
    ca_654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_308_inst_ack_1, ack => maxPool4_CP_563_elements(29)); -- 
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	13 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 call_stmt_293_to_assign_stmt_792/slice_312_sample_start_
      -- CP-element group 30: 	 call_stmt_293_to_assign_stmt_792/slice_312_Sample/rr
      -- CP-element group 30: 	 call_stmt_293_to_assign_stmt_792/slice_312_Sample/$entry
      -- 
    rr_662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(30), ack => slice_312_inst_req_0); -- 
    maxPool4_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(13) & maxPool4_CP_563_elements(32);
      gj_maxPool4_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: 	164 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 call_stmt_293_to_assign_stmt_792/slice_312_Update/cr
      -- CP-element group 31: 	 call_stmt_293_to_assign_stmt_792/slice_312_Update/$entry
      -- CP-element group 31: 	 call_stmt_293_to_assign_stmt_792/slice_312_update_start_
      -- 
    cr_667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(31), ack => slice_312_inst_req_1); -- 
    maxPool4_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(33) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	11 
    -- CP-element group 32: 	30 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 call_stmt_293_to_assign_stmt_792/slice_312_sample_completed_
      -- CP-element group 32: 	 call_stmt_293_to_assign_stmt_792/slice_312_Sample/ra
      -- CP-element group 32: 	 call_stmt_293_to_assign_stmt_792/slice_312_Sample/$exit
      -- 
    ra_663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_312_inst_ack_0, ack => maxPool4_CP_563_elements(32)); -- 
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	162 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 call_stmt_293_to_assign_stmt_792/slice_312_Update/$exit
      -- CP-element group 33: 	 call_stmt_293_to_assign_stmt_792/slice_312_Update/ca
      -- CP-element group 33: 	 call_stmt_293_to_assign_stmt_792/slice_312_update_completed_
      -- 
    ca_668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_312_inst_ack_1, ack => maxPool4_CP_563_elements(33)); -- 
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 call_stmt_293_to_assign_stmt_792/slice_316_Sample/rr
      -- CP-element group 34: 	 call_stmt_293_to_assign_stmt_792/slice_316_Sample/$entry
      -- CP-element group 34: 	 call_stmt_293_to_assign_stmt_792/slice_316_sample_start_
      -- 
    rr_676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(34), ack => slice_316_inst_req_0); -- 
    maxPool4_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(13) & maxPool4_CP_563_elements(36);
      gj_maxPool4_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	37 
    -- CP-element group 35: 	164 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 call_stmt_293_to_assign_stmt_792/slice_316_update_start_
      -- CP-element group 35: 	 call_stmt_293_to_assign_stmt_792/slice_316_Update/cr
      -- CP-element group 35: 	 call_stmt_293_to_assign_stmt_792/slice_316_Update/$entry
      -- 
    cr_681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(35), ack => slice_316_inst_req_1); -- 
    maxPool4_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(37) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: 	34 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 call_stmt_293_to_assign_stmt_792/slice_316_sample_completed_
      -- CP-element group 36: 	 call_stmt_293_to_assign_stmt_792/slice_316_Sample/ra
      -- CP-element group 36: 	 call_stmt_293_to_assign_stmt_792/slice_316_Sample/$exit
      -- 
    ra_677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_316_inst_ack_0, ack => maxPool4_CP_563_elements(36)); -- 
    -- CP-element group 37:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	162 
    -- CP-element group 37: marked-successors 
    -- CP-element group 37: 	35 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 call_stmt_293_to_assign_stmt_792/slice_316_update_completed_
      -- CP-element group 37: 	 call_stmt_293_to_assign_stmt_792/slice_316_Update/ca
      -- CP-element group 37: 	 call_stmt_293_to_assign_stmt_792/slice_316_Update/$exit
      -- 
    ca_682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_316_inst_ack_1, ack => maxPool4_CP_563_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	40 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 call_stmt_293_to_assign_stmt_792/slice_320_sample_start_
      -- CP-element group 38: 	 call_stmt_293_to_assign_stmt_792/slice_320_Sample/rr
      -- CP-element group 38: 	 call_stmt_293_to_assign_stmt_792/slice_320_Sample/$entry
      -- 
    rr_690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(38), ack => slice_320_inst_req_0); -- 
    maxPool4_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(13) & maxPool4_CP_563_elements(40);
      gj_maxPool4_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: 	164 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 call_stmt_293_to_assign_stmt_792/slice_320_Update/$entry
      -- CP-element group 39: 	 call_stmt_293_to_assign_stmt_792/slice_320_Update/cr
      -- CP-element group 39: 	 call_stmt_293_to_assign_stmt_792/slice_320_update_start_
      -- 
    cr_695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(39), ack => slice_320_inst_req_1); -- 
    maxPool4_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(41) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: 	11 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 call_stmt_293_to_assign_stmt_792/slice_320_sample_completed_
      -- CP-element group 40: 	 call_stmt_293_to_assign_stmt_792/slice_320_Sample/ra
      -- CP-element group 40: 	 call_stmt_293_to_assign_stmt_792/slice_320_Sample/$exit
      -- 
    ra_691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_320_inst_ack_0, ack => maxPool4_CP_563_elements(40)); -- 
    -- CP-element group 41:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	162 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	39 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 call_stmt_293_to_assign_stmt_792/slice_320_Update/$exit
      -- CP-element group 41: 	 call_stmt_293_to_assign_stmt_792/slice_320_update_completed_
      -- CP-element group 41: 	 call_stmt_293_to_assign_stmt_792/slice_320_Update/ca
      -- 
    ca_696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_320_inst_ack_1, ack => maxPool4_CP_563_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	13 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 call_stmt_293_to_assign_stmt_792/slice_324_sample_start_
      -- CP-element group 42: 	 call_stmt_293_to_assign_stmt_792/slice_324_Sample/rr
      -- CP-element group 42: 	 call_stmt_293_to_assign_stmt_792/slice_324_Sample/$entry
      -- 
    rr_704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(42), ack => slice_324_inst_req_0); -- 
    maxPool4_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(13) & maxPool4_CP_563_elements(44);
      gj_maxPool4_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	45 
    -- CP-element group 43: 	164 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 call_stmt_293_to_assign_stmt_792/slice_324_Update/cr
      -- CP-element group 43: 	 call_stmt_293_to_assign_stmt_792/slice_324_Update/$entry
      -- CP-element group 43: 	 call_stmt_293_to_assign_stmt_792/slice_324_update_start_
      -- 
    cr_709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(43), ack => slice_324_inst_req_1); -- 
    maxPool4_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(45) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: 	11 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 call_stmt_293_to_assign_stmt_792/slice_324_sample_completed_
      -- CP-element group 44: 	 call_stmt_293_to_assign_stmt_792/slice_324_Sample/ra
      -- CP-element group 44: 	 call_stmt_293_to_assign_stmt_792/slice_324_Sample/$exit
      -- 
    ra_705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_324_inst_ack_0, ack => maxPool4_CP_563_elements(44)); -- 
    -- CP-element group 45:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	162 
    -- CP-element group 45: marked-successors 
    -- CP-element group 45: 	43 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 call_stmt_293_to_assign_stmt_792/slice_324_Update/ca
      -- CP-element group 45: 	 call_stmt_293_to_assign_stmt_792/slice_324_Update/$exit
      -- CP-element group 45: 	 call_stmt_293_to_assign_stmt_792/slice_324_update_completed_
      -- 
    ca_710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_324_inst_ack_1, ack => maxPool4_CP_563_elements(45)); -- 
    -- CP-element group 46:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	13 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	48 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 call_stmt_293_to_assign_stmt_792/slice_328_Sample/rr
      -- CP-element group 46: 	 call_stmt_293_to_assign_stmt_792/slice_328_Sample/$entry
      -- CP-element group 46: 	 call_stmt_293_to_assign_stmt_792/slice_328_sample_start_
      -- 
    rr_718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(46), ack => slice_328_inst_req_0); -- 
    maxPool4_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(13) & maxPool4_CP_563_elements(48);
      gj_maxPool4_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	49 
    -- CP-element group 47: 	164 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 call_stmt_293_to_assign_stmt_792/slice_328_Update/cr
      -- CP-element group 47: 	 call_stmt_293_to_assign_stmt_792/slice_328_Update/$entry
      -- CP-element group 47: 	 call_stmt_293_to_assign_stmt_792/slice_328_update_start_
      -- 
    cr_723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(47), ack => slice_328_inst_req_1); -- 
    maxPool4_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(49) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: marked-successors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: 	11 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 call_stmt_293_to_assign_stmt_792/slice_328_Sample/ra
      -- CP-element group 48: 	 call_stmt_293_to_assign_stmt_792/slice_328_Sample/$exit
      -- CP-element group 48: 	 call_stmt_293_to_assign_stmt_792/slice_328_sample_completed_
      -- 
    ra_719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_328_inst_ack_0, ack => maxPool4_CP_563_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	162 
    -- CP-element group 49: marked-successors 
    -- CP-element group 49: 	47 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 call_stmt_293_to_assign_stmt_792/slice_328_Update/ca
      -- CP-element group 49: 	 call_stmt_293_to_assign_stmt_792/slice_328_Update/$exit
      -- CP-element group 49: 	 call_stmt_293_to_assign_stmt_792/slice_328_update_completed_
      -- 
    ca_724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_328_inst_ack_1, ack => maxPool4_CP_563_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	13 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	52 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 call_stmt_293_to_assign_stmt_792/slice_332_sample_start_
      -- CP-element group 50: 	 call_stmt_293_to_assign_stmt_792/slice_332_Sample/rr
      -- CP-element group 50: 	 call_stmt_293_to_assign_stmt_792/slice_332_Sample/$entry
      -- 
    rr_732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(50), ack => slice_332_inst_req_0); -- 
    maxPool4_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(13) & maxPool4_CP_563_elements(52);
      gj_maxPool4_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	53 
    -- CP-element group 51: 	164 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 call_stmt_293_to_assign_stmt_792/slice_332_Update/cr
      -- CP-element group 51: 	 call_stmt_293_to_assign_stmt_792/slice_332_Update/$entry
      -- CP-element group 51: 	 call_stmt_293_to_assign_stmt_792/slice_332_update_start_
      -- 
    cr_737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(51), ack => slice_332_inst_req_1); -- 
    maxPool4_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(53) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: 	11 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 call_stmt_293_to_assign_stmt_792/slice_332_Sample/ra
      -- CP-element group 52: 	 call_stmt_293_to_assign_stmt_792/slice_332_sample_completed_
      -- CP-element group 52: 	 call_stmt_293_to_assign_stmt_792/slice_332_Sample/$exit
      -- 
    ra_733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_332_inst_ack_0, ack => maxPool4_CP_563_elements(52)); -- 
    -- CP-element group 53:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	162 
    -- CP-element group 53: marked-successors 
    -- CP-element group 53: 	51 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 call_stmt_293_to_assign_stmt_792/slice_332_Update/$exit
      -- CP-element group 53: 	 call_stmt_293_to_assign_stmt_792/slice_332_update_completed_
      -- CP-element group 53: 	 call_stmt_293_to_assign_stmt_792/slice_332_Update/ca
      -- 
    ca_738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_332_inst_ack_1, ack => maxPool4_CP_563_elements(53)); -- 
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	13 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	56 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 call_stmt_293_to_assign_stmt_792/slice_336_Sample/rr
      -- CP-element group 54: 	 call_stmt_293_to_assign_stmt_792/slice_336_Sample/$entry
      -- CP-element group 54: 	 call_stmt_293_to_assign_stmt_792/slice_336_sample_start_
      -- 
    rr_746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(54), ack => slice_336_inst_req_0); -- 
    maxPool4_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(13) & maxPool4_CP_563_elements(56);
      gj_maxPool4_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	57 
    -- CP-element group 55: 	164 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 call_stmt_293_to_assign_stmt_792/slice_336_Update/$entry
      -- CP-element group 55: 	 call_stmt_293_to_assign_stmt_792/slice_336_update_start_
      -- CP-element group 55: 	 call_stmt_293_to_assign_stmt_792/slice_336_Update/cr
      -- 
    cr_751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(55), ack => slice_336_inst_req_1); -- 
    maxPool4_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(57) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: 	11 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 call_stmt_293_to_assign_stmt_792/slice_336_Sample/ra
      -- CP-element group 56: 	 call_stmt_293_to_assign_stmt_792/slice_336_sample_completed_
      -- CP-element group 56: 	 call_stmt_293_to_assign_stmt_792/slice_336_Sample/$exit
      -- 
    ra_747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_336_inst_ack_0, ack => maxPool4_CP_563_elements(56)); -- 
    -- CP-element group 57:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	162 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	55 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 call_stmt_293_to_assign_stmt_792/slice_336_update_completed_
      -- CP-element group 57: 	 call_stmt_293_to_assign_stmt_792/slice_336_Update/$exit
      -- CP-element group 57: 	 call_stmt_293_to_assign_stmt_792/slice_336_Update/ca
      -- 
    ca_752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_336_inst_ack_1, ack => maxPool4_CP_563_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	17 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 call_stmt_293_to_assign_stmt_792/slice_340_Sample/$entry
      -- CP-element group 58: 	 call_stmt_293_to_assign_stmt_792/slice_340_sample_start_
      -- CP-element group 58: 	 call_stmt_293_to_assign_stmt_792/slice_340_Sample/rr
      -- 
    rr_760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(58), ack => slice_340_inst_req_0); -- 
    maxPool4_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(17) & maxPool4_CP_563_elements(60);
      gj_maxPool4_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: 	164 
    -- CP-element group 59: 	168 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 call_stmt_293_to_assign_stmt_792/slice_340_update_start_
      -- CP-element group 59: 	 call_stmt_293_to_assign_stmt_792/slice_340_Update/cr
      -- CP-element group 59: 	 call_stmt_293_to_assign_stmt_792/slice_340_Update/$entry
      -- 
    cr_765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(59), ack => slice_340_inst_req_1); -- 
    maxPool4_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(61) & maxPool4_CP_563_elements(164) & maxPool4_CP_563_elements(168);
      gj_maxPool4_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: 	15 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 call_stmt_293_to_assign_stmt_792/slice_340_sample_completed_
      -- CP-element group 60: 	 call_stmt_293_to_assign_stmt_792/slice_340_Sample/$exit
      -- CP-element group 60: 	 call_stmt_293_to_assign_stmt_792/slice_340_Sample/ra
      -- 
    ra_761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_340_inst_ack_0, ack => maxPool4_CP_563_elements(60)); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	162 
    -- CP-element group 61: 	166 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 call_stmt_293_to_assign_stmt_792/slice_340_update_completed_
      -- CP-element group 61: 	 call_stmt_293_to_assign_stmt_792/slice_340_Update/ca
      -- CP-element group 61: 	 call_stmt_293_to_assign_stmt_792/slice_340_Update/$exit
      -- 
    ca_766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_340_inst_ack_1, ack => maxPool4_CP_563_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	17 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 call_stmt_293_to_assign_stmt_792/slice_344_Sample/rr
      -- CP-element group 62: 	 call_stmt_293_to_assign_stmt_792/slice_344_sample_start_
      -- CP-element group 62: 	 call_stmt_293_to_assign_stmt_792/slice_344_Sample/$entry
      -- 
    rr_774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(62), ack => slice_344_inst_req_0); -- 
    maxPool4_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(17) & maxPool4_CP_563_elements(64);
      gj_maxPool4_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: 	164 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 call_stmt_293_to_assign_stmt_792/slice_344_Update/cr
      -- CP-element group 63: 	 call_stmt_293_to_assign_stmt_792/slice_344_update_start_
      -- CP-element group 63: 	 call_stmt_293_to_assign_stmt_792/slice_344_Update/$entry
      -- 
    cr_779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(63), ack => slice_344_inst_req_1); -- 
    maxPool4_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(65) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: 	15 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 call_stmt_293_to_assign_stmt_792/slice_344_Sample/ra
      -- CP-element group 64: 	 call_stmt_293_to_assign_stmt_792/slice_344_sample_completed_
      -- CP-element group 64: 	 call_stmt_293_to_assign_stmt_792/slice_344_Sample/$exit
      -- 
    ra_775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_344_inst_ack_0, ack => maxPool4_CP_563_elements(64)); -- 
    -- CP-element group 65:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	162 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	63 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 call_stmt_293_to_assign_stmt_792/slice_344_Update/ca
      -- CP-element group 65: 	 call_stmt_293_to_assign_stmt_792/slice_344_Update/$exit
      -- CP-element group 65: 	 call_stmt_293_to_assign_stmt_792/slice_344_update_completed_
      -- 
    ca_780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_344_inst_ack_1, ack => maxPool4_CP_563_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	17 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	68 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 call_stmt_293_to_assign_stmt_792/slice_348_Sample/rr
      -- CP-element group 66: 	 call_stmt_293_to_assign_stmt_792/slice_348_sample_start_
      -- CP-element group 66: 	 call_stmt_293_to_assign_stmt_792/slice_348_Sample/$entry
      -- 
    rr_788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(66), ack => slice_348_inst_req_0); -- 
    maxPool4_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(17) & maxPool4_CP_563_elements(68);
      gj_maxPool4_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: 	164 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 call_stmt_293_to_assign_stmt_792/slice_348_Update/$entry
      -- CP-element group 67: 	 call_stmt_293_to_assign_stmt_792/slice_348_update_start_
      -- CP-element group 67: 	 call_stmt_293_to_assign_stmt_792/slice_348_Update/cr
      -- 
    cr_793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(67), ack => slice_348_inst_req_1); -- 
    maxPool4_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(69) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: 	15 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 call_stmt_293_to_assign_stmt_792/slice_348_Sample/ra
      -- CP-element group 68: 	 call_stmt_293_to_assign_stmt_792/slice_348_sample_completed_
      -- CP-element group 68: 	 call_stmt_293_to_assign_stmt_792/slice_348_Sample/$exit
      -- 
    ra_789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_348_inst_ack_0, ack => maxPool4_CP_563_elements(68)); -- 
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	162 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	67 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 call_stmt_293_to_assign_stmt_792/slice_348_update_completed_
      -- CP-element group 69: 	 call_stmt_293_to_assign_stmt_792/slice_348_Update/$exit
      -- CP-element group 69: 	 call_stmt_293_to_assign_stmt_792/slice_348_Update/ca
      -- 
    ca_794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_348_inst_ack_1, ack => maxPool4_CP_563_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	17 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	72 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 call_stmt_293_to_assign_stmt_792/slice_352_Sample/$entry
      -- CP-element group 70: 	 call_stmt_293_to_assign_stmt_792/slice_352_Sample/rr
      -- CP-element group 70: 	 call_stmt_293_to_assign_stmt_792/slice_352_sample_start_
      -- 
    rr_802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(70), ack => slice_352_inst_req_0); -- 
    maxPool4_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(17) & maxPool4_CP_563_elements(72);
      gj_maxPool4_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: 	164 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 call_stmt_293_to_assign_stmt_792/slice_352_update_start_
      -- CP-element group 71: 	 call_stmt_293_to_assign_stmt_792/slice_352_Update/cr
      -- CP-element group 71: 	 call_stmt_293_to_assign_stmt_792/slice_352_Update/$entry
      -- 
    cr_807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(71), ack => slice_352_inst_req_1); -- 
    maxPool4_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(73) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: 	15 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 call_stmt_293_to_assign_stmt_792/slice_352_Sample/$exit
      -- CP-element group 72: 	 call_stmt_293_to_assign_stmt_792/slice_352_sample_completed_
      -- CP-element group 72: 	 call_stmt_293_to_assign_stmt_792/slice_352_Sample/ra
      -- 
    ra_803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_352_inst_ack_0, ack => maxPool4_CP_563_elements(72)); -- 
    -- CP-element group 73:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	162 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	71 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 call_stmt_293_to_assign_stmt_792/slice_352_update_completed_
      -- CP-element group 73: 	 call_stmt_293_to_assign_stmt_792/slice_352_Update/$exit
      -- CP-element group 73: 	 call_stmt_293_to_assign_stmt_792/slice_352_Update/ca
      -- 
    ca_808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_352_inst_ack_1, ack => maxPool4_CP_563_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	17 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 call_stmt_293_to_assign_stmt_792/slice_356_Sample/$entry
      -- CP-element group 74: 	 call_stmt_293_to_assign_stmt_792/slice_356_Sample/rr
      -- CP-element group 74: 	 call_stmt_293_to_assign_stmt_792/slice_356_sample_start_
      -- 
    rr_816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(74), ack => slice_356_inst_req_0); -- 
    maxPool4_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(17) & maxPool4_CP_563_elements(76);
      gj_maxPool4_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: 	164 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 call_stmt_293_to_assign_stmt_792/slice_356_Update/cr
      -- CP-element group 75: 	 call_stmt_293_to_assign_stmt_792/slice_356_update_start_
      -- CP-element group 75: 	 call_stmt_293_to_assign_stmt_792/slice_356_Update/$entry
      -- 
    cr_821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(75), ack => slice_356_inst_req_1); -- 
    maxPool4_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(77) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	15 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 call_stmt_293_to_assign_stmt_792/slice_356_Sample/$exit
      -- CP-element group 76: 	 call_stmt_293_to_assign_stmt_792/slice_356_sample_completed_
      -- CP-element group 76: 	 call_stmt_293_to_assign_stmt_792/slice_356_Sample/ra
      -- 
    ra_817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_356_inst_ack_0, ack => maxPool4_CP_563_elements(76)); -- 
    -- CP-element group 77:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	162 
    -- CP-element group 77: marked-successors 
    -- CP-element group 77: 	75 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 call_stmt_293_to_assign_stmt_792/slice_356_Update/ca
      -- CP-element group 77: 	 call_stmt_293_to_assign_stmt_792/slice_356_update_completed_
      -- CP-element group 77: 	 call_stmt_293_to_assign_stmt_792/slice_356_Update/$exit
      -- 
    ca_822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_356_inst_ack_1, ack => maxPool4_CP_563_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	17 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	80 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 call_stmt_293_to_assign_stmt_792/slice_360_sample_start_
      -- CP-element group 78: 	 call_stmt_293_to_assign_stmt_792/slice_360_Sample/$entry
      -- CP-element group 78: 	 call_stmt_293_to_assign_stmt_792/slice_360_Sample/rr
      -- 
    rr_830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(78), ack => slice_360_inst_req_0); -- 
    maxPool4_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(17) & maxPool4_CP_563_elements(80);
      gj_maxPool4_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	81 
    -- CP-element group 79: 	164 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 call_stmt_293_to_assign_stmt_792/slice_360_update_start_
      -- CP-element group 79: 	 call_stmt_293_to_assign_stmt_792/slice_360_Update/$entry
      -- CP-element group 79: 	 call_stmt_293_to_assign_stmt_792/slice_360_Update/cr
      -- 
    cr_835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(79), ack => slice_360_inst_req_1); -- 
    maxPool4_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(81) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	15 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 call_stmt_293_to_assign_stmt_792/slice_360_sample_completed_
      -- CP-element group 80: 	 call_stmt_293_to_assign_stmt_792/slice_360_Sample/$exit
      -- CP-element group 80: 	 call_stmt_293_to_assign_stmt_792/slice_360_Sample/ra
      -- 
    ra_831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_360_inst_ack_0, ack => maxPool4_CP_563_elements(80)); -- 
    -- CP-element group 81:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	162 
    -- CP-element group 81: marked-successors 
    -- CP-element group 81: 	79 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 call_stmt_293_to_assign_stmt_792/slice_360_update_completed_
      -- CP-element group 81: 	 call_stmt_293_to_assign_stmt_792/slice_360_Update/$exit
      -- CP-element group 81: 	 call_stmt_293_to_assign_stmt_792/slice_360_Update/ca
      -- 
    ca_836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_360_inst_ack_1, ack => maxPool4_CP_563_elements(81)); -- 
    -- CP-element group 82:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	17 
    -- CP-element group 82: marked-predecessors 
    -- CP-element group 82: 	84 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 call_stmt_293_to_assign_stmt_792/slice_364_sample_start_
      -- CP-element group 82: 	 call_stmt_293_to_assign_stmt_792/slice_364_Sample/$entry
      -- CP-element group 82: 	 call_stmt_293_to_assign_stmt_792/slice_364_Sample/rr
      -- 
    rr_844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(82), ack => slice_364_inst_req_0); -- 
    maxPool4_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(17) & maxPool4_CP_563_elements(84);
      gj_maxPool4_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: 	164 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 call_stmt_293_to_assign_stmt_792/slice_364_Update/$entry
      -- CP-element group 83: 	 call_stmt_293_to_assign_stmt_792/slice_364_update_start_
      -- CP-element group 83: 	 call_stmt_293_to_assign_stmt_792/slice_364_Update/cr
      -- 
    cr_849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(83), ack => slice_364_inst_req_1); -- 
    maxPool4_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(85) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: marked-successors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	15 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 call_stmt_293_to_assign_stmt_792/slice_364_sample_completed_
      -- CP-element group 84: 	 call_stmt_293_to_assign_stmt_792/slice_364_Sample/$exit
      -- CP-element group 84: 	 call_stmt_293_to_assign_stmt_792/slice_364_Sample/ra
      -- 
    ra_845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_364_inst_ack_0, ack => maxPool4_CP_563_elements(84)); -- 
    -- CP-element group 85:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	162 
    -- CP-element group 85: marked-successors 
    -- CP-element group 85: 	83 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 call_stmt_293_to_assign_stmt_792/slice_364_update_completed_
      -- CP-element group 85: 	 call_stmt_293_to_assign_stmt_792/slice_364_Update/$exit
      -- CP-element group 85: 	 call_stmt_293_to_assign_stmt_792/slice_364_Update/ca
      -- 
    ca_850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_364_inst_ack_1, ack => maxPool4_CP_563_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	17 
    -- CP-element group 86: marked-predecessors 
    -- CP-element group 86: 	88 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 call_stmt_293_to_assign_stmt_792/slice_368_sample_start_
      -- CP-element group 86: 	 call_stmt_293_to_assign_stmt_792/slice_368_Sample/$entry
      -- CP-element group 86: 	 call_stmt_293_to_assign_stmt_792/slice_368_Sample/rr
      -- 
    rr_858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(86), ack => slice_368_inst_req_0); -- 
    maxPool4_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(17) & maxPool4_CP_563_elements(88);
      gj_maxPool4_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: marked-predecessors 
    -- CP-element group 87: 	89 
    -- CP-element group 87: 	164 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 call_stmt_293_to_assign_stmt_792/slice_368_update_start_
      -- CP-element group 87: 	 call_stmt_293_to_assign_stmt_792/slice_368_Update/$entry
      -- CP-element group 87: 	 call_stmt_293_to_assign_stmt_792/slice_368_Update/cr
      -- 
    cr_863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(87), ack => slice_368_inst_req_1); -- 
    maxPool4_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(89) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: marked-successors 
    -- CP-element group 88: 	15 
    -- CP-element group 88: 	86 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 call_stmt_293_to_assign_stmt_792/slice_368_sample_completed_
      -- CP-element group 88: 	 call_stmt_293_to_assign_stmt_792/slice_368_Sample/$exit
      -- CP-element group 88: 	 call_stmt_293_to_assign_stmt_792/slice_368_Sample/ra
      -- 
    ra_859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_368_inst_ack_0, ack => maxPool4_CP_563_elements(88)); -- 
    -- CP-element group 89:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	162 
    -- CP-element group 89: marked-successors 
    -- CP-element group 89: 	87 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 call_stmt_293_to_assign_stmt_792/slice_368_update_completed_
      -- CP-element group 89: 	 call_stmt_293_to_assign_stmt_792/slice_368_Update/$exit
      -- CP-element group 89: 	 call_stmt_293_to_assign_stmt_792/slice_368_Update/ca
      -- 
    ca_864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_368_inst_ack_1, ack => maxPool4_CP_563_elements(89)); -- 
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	21 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	92 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 call_stmt_293_to_assign_stmt_792/slice_372_sample_start_
      -- CP-element group 90: 	 call_stmt_293_to_assign_stmt_792/slice_372_Sample/$entry
      -- CP-element group 90: 	 call_stmt_293_to_assign_stmt_792/slice_372_Sample/rr
      -- 
    rr_872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(90), ack => slice_372_inst_req_0); -- 
    maxPool4_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(21) & maxPool4_CP_563_elements(92);
      gj_maxPool4_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: marked-predecessors 
    -- CP-element group 91: 	93 
    -- CP-element group 91: 	164 
    -- CP-element group 91: 	168 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 call_stmt_293_to_assign_stmt_792/slice_372_update_start_
      -- CP-element group 91: 	 call_stmt_293_to_assign_stmt_792/slice_372_Update/$entry
      -- CP-element group 91: 	 call_stmt_293_to_assign_stmt_792/slice_372_Update/cr
      -- 
    cr_877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(91), ack => slice_372_inst_req_1); -- 
    maxPool4_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(93) & maxPool4_CP_563_elements(164) & maxPool4_CP_563_elements(168);
      gj_maxPool4_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: marked-successors 
    -- CP-element group 92: 	19 
    -- CP-element group 92: 	90 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 call_stmt_293_to_assign_stmt_792/slice_372_sample_completed_
      -- CP-element group 92: 	 call_stmt_293_to_assign_stmt_792/slice_372_Sample/$exit
      -- CP-element group 92: 	 call_stmt_293_to_assign_stmt_792/slice_372_Sample/ra
      -- 
    ra_873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_372_inst_ack_0, ack => maxPool4_CP_563_elements(92)); -- 
    -- CP-element group 93:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	162 
    -- CP-element group 93: 	166 
    -- CP-element group 93: marked-successors 
    -- CP-element group 93: 	91 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 call_stmt_293_to_assign_stmt_792/slice_372_update_completed_
      -- CP-element group 93: 	 call_stmt_293_to_assign_stmt_792/slice_372_Update/$exit
      -- CP-element group 93: 	 call_stmt_293_to_assign_stmt_792/slice_372_Update/ca
      -- 
    ca_878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_372_inst_ack_1, ack => maxPool4_CP_563_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	21 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	96 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 call_stmt_293_to_assign_stmt_792/slice_376_sample_start_
      -- CP-element group 94: 	 call_stmt_293_to_assign_stmt_792/slice_376_Sample/$entry
      -- CP-element group 94: 	 call_stmt_293_to_assign_stmt_792/slice_376_Sample/rr
      -- 
    rr_886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(94), ack => slice_376_inst_req_0); -- 
    maxPool4_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(21) & maxPool4_CP_563_elements(96);
      gj_maxPool4_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	97 
    -- CP-element group 95: 	164 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 call_stmt_293_to_assign_stmt_792/slice_376_update_start_
      -- CP-element group 95: 	 call_stmt_293_to_assign_stmt_792/slice_376_Update/$entry
      -- CP-element group 95: 	 call_stmt_293_to_assign_stmt_792/slice_376_Update/cr
      -- 
    cr_891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(95), ack => slice_376_inst_req_1); -- 
    maxPool4_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(97) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	19 
    -- CP-element group 96: 	94 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 call_stmt_293_to_assign_stmt_792/slice_376_sample_completed_
      -- CP-element group 96: 	 call_stmt_293_to_assign_stmt_792/slice_376_Sample/$exit
      -- CP-element group 96: 	 call_stmt_293_to_assign_stmt_792/slice_376_Sample/ra
      -- 
    ra_887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_376_inst_ack_0, ack => maxPool4_CP_563_elements(96)); -- 
    -- CP-element group 97:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	162 
    -- CP-element group 97: marked-successors 
    -- CP-element group 97: 	95 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 call_stmt_293_to_assign_stmt_792/slice_376_update_completed_
      -- CP-element group 97: 	 call_stmt_293_to_assign_stmt_792/slice_376_Update/$exit
      -- CP-element group 97: 	 call_stmt_293_to_assign_stmt_792/slice_376_Update/ca
      -- 
    ca_892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_376_inst_ack_1, ack => maxPool4_CP_563_elements(97)); -- 
    -- CP-element group 98:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	21 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	100 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 call_stmt_293_to_assign_stmt_792/slice_380_sample_start_
      -- CP-element group 98: 	 call_stmt_293_to_assign_stmt_792/slice_380_Sample/$entry
      -- CP-element group 98: 	 call_stmt_293_to_assign_stmt_792/slice_380_Sample/rr
      -- 
    rr_900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(98), ack => slice_380_inst_req_0); -- 
    maxPool4_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(21) & maxPool4_CP_563_elements(100);
      gj_maxPool4_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: marked-predecessors 
    -- CP-element group 99: 	101 
    -- CP-element group 99: 	164 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 call_stmt_293_to_assign_stmt_792/slice_380_update_start_
      -- CP-element group 99: 	 call_stmt_293_to_assign_stmt_792/slice_380_Update/$entry
      -- CP-element group 99: 	 call_stmt_293_to_assign_stmt_792/slice_380_Update/cr
      -- 
    cr_905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(99), ack => slice_380_inst_req_1); -- 
    maxPool4_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(101) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_99 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: successors 
    -- CP-element group 100: marked-successors 
    -- CP-element group 100: 	19 
    -- CP-element group 100: 	98 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 call_stmt_293_to_assign_stmt_792/slice_380_sample_completed_
      -- CP-element group 100: 	 call_stmt_293_to_assign_stmt_792/slice_380_Sample/$exit
      -- CP-element group 100: 	 call_stmt_293_to_assign_stmt_792/slice_380_Sample/ra
      -- 
    ra_901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_380_inst_ack_0, ack => maxPool4_CP_563_elements(100)); -- 
    -- CP-element group 101:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	162 
    -- CP-element group 101: marked-successors 
    -- CP-element group 101: 	99 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 call_stmt_293_to_assign_stmt_792/slice_380_update_completed_
      -- CP-element group 101: 	 call_stmt_293_to_assign_stmt_792/slice_380_Update/$exit
      -- CP-element group 101: 	 call_stmt_293_to_assign_stmt_792/slice_380_Update/ca
      -- 
    ca_906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_380_inst_ack_1, ack => maxPool4_CP_563_elements(101)); -- 
    -- CP-element group 102:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	21 
    -- CP-element group 102: marked-predecessors 
    -- CP-element group 102: 	104 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 call_stmt_293_to_assign_stmt_792/slice_384_sample_start_
      -- CP-element group 102: 	 call_stmt_293_to_assign_stmt_792/slice_384_Sample/$entry
      -- CP-element group 102: 	 call_stmt_293_to_assign_stmt_792/slice_384_Sample/rr
      -- 
    rr_914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(102), ack => slice_384_inst_req_0); -- 
    maxPool4_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(21) & maxPool4_CP_563_elements(104);
      gj_maxPool4_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: marked-predecessors 
    -- CP-element group 103: 	105 
    -- CP-element group 103: 	164 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 call_stmt_293_to_assign_stmt_792/slice_384_update_start_
      -- CP-element group 103: 	 call_stmt_293_to_assign_stmt_792/slice_384_Update/$entry
      -- CP-element group 103: 	 call_stmt_293_to_assign_stmt_792/slice_384_Update/cr
      -- 
    cr_919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(103), ack => slice_384_inst_req_1); -- 
    maxPool4_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(105) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104: marked-successors 
    -- CP-element group 104: 	19 
    -- CP-element group 104: 	102 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 call_stmt_293_to_assign_stmt_792/slice_384_sample_completed_
      -- CP-element group 104: 	 call_stmt_293_to_assign_stmt_792/slice_384_Sample/$exit
      -- CP-element group 104: 	 call_stmt_293_to_assign_stmt_792/slice_384_Sample/ra
      -- 
    ra_915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_384_inst_ack_0, ack => maxPool4_CP_563_elements(104)); -- 
    -- CP-element group 105:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	162 
    -- CP-element group 105: marked-successors 
    -- CP-element group 105: 	103 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 call_stmt_293_to_assign_stmt_792/slice_384_update_completed_
      -- CP-element group 105: 	 call_stmt_293_to_assign_stmt_792/slice_384_Update/$exit
      -- CP-element group 105: 	 call_stmt_293_to_assign_stmt_792/slice_384_Update/ca
      -- 
    ca_920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_384_inst_ack_1, ack => maxPool4_CP_563_elements(105)); -- 
    -- CP-element group 106:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	21 
    -- CP-element group 106: marked-predecessors 
    -- CP-element group 106: 	108 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 call_stmt_293_to_assign_stmt_792/slice_388_sample_start_
      -- CP-element group 106: 	 call_stmt_293_to_assign_stmt_792/slice_388_Sample/$entry
      -- CP-element group 106: 	 call_stmt_293_to_assign_stmt_792/slice_388_Sample/rr
      -- 
    rr_928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(106), ack => slice_388_inst_req_0); -- 
    maxPool4_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(21) & maxPool4_CP_563_elements(108);
      gj_maxPool4_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: marked-predecessors 
    -- CP-element group 107: 	109 
    -- CP-element group 107: 	164 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 call_stmt_293_to_assign_stmt_792/slice_388_update_start_
      -- CP-element group 107: 	 call_stmt_293_to_assign_stmt_792/slice_388_Update/$entry
      -- CP-element group 107: 	 call_stmt_293_to_assign_stmt_792/slice_388_Update/cr
      -- 
    cr_933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(107), ack => slice_388_inst_req_1); -- 
    maxPool4_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(109) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108: marked-successors 
    -- CP-element group 108: 	19 
    -- CP-element group 108: 	106 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 call_stmt_293_to_assign_stmt_792/slice_388_sample_completed_
      -- CP-element group 108: 	 call_stmt_293_to_assign_stmt_792/slice_388_Sample/$exit
      -- CP-element group 108: 	 call_stmt_293_to_assign_stmt_792/slice_388_Sample/ra
      -- 
    ra_929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_388_inst_ack_0, ack => maxPool4_CP_563_elements(108)); -- 
    -- CP-element group 109:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	162 
    -- CP-element group 109: marked-successors 
    -- CP-element group 109: 	107 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 call_stmt_293_to_assign_stmt_792/slice_388_update_completed_
      -- CP-element group 109: 	 call_stmt_293_to_assign_stmt_792/slice_388_Update/$exit
      -- CP-element group 109: 	 call_stmt_293_to_assign_stmt_792/slice_388_Update/ca
      -- 
    ca_934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_388_inst_ack_1, ack => maxPool4_CP_563_elements(109)); -- 
    -- CP-element group 110:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	21 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	112 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 call_stmt_293_to_assign_stmt_792/slice_392_sample_start_
      -- CP-element group 110: 	 call_stmt_293_to_assign_stmt_792/slice_392_Sample/$entry
      -- CP-element group 110: 	 call_stmt_293_to_assign_stmt_792/slice_392_Sample/rr
      -- 
    rr_942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(110), ack => slice_392_inst_req_0); -- 
    maxPool4_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(21) & maxPool4_CP_563_elements(112);
      gj_maxPool4_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: marked-predecessors 
    -- CP-element group 111: 	113 
    -- CP-element group 111: 	164 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 call_stmt_293_to_assign_stmt_792/slice_392_update_start_
      -- CP-element group 111: 	 call_stmt_293_to_assign_stmt_792/slice_392_Update/$entry
      -- CP-element group 111: 	 call_stmt_293_to_assign_stmt_792/slice_392_Update/cr
      -- 
    cr_947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(111), ack => slice_392_inst_req_1); -- 
    maxPool4_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(113) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: marked-successors 
    -- CP-element group 112: 	19 
    -- CP-element group 112: 	110 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 call_stmt_293_to_assign_stmt_792/slice_392_sample_completed_
      -- CP-element group 112: 	 call_stmt_293_to_assign_stmt_792/slice_392_Sample/$exit
      -- CP-element group 112: 	 call_stmt_293_to_assign_stmt_792/slice_392_Sample/ra
      -- 
    ra_943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_392_inst_ack_0, ack => maxPool4_CP_563_elements(112)); -- 
    -- CP-element group 113:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	162 
    -- CP-element group 113: marked-successors 
    -- CP-element group 113: 	111 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 call_stmt_293_to_assign_stmt_792/slice_392_update_completed_
      -- CP-element group 113: 	 call_stmt_293_to_assign_stmt_792/slice_392_Update/$exit
      -- CP-element group 113: 	 call_stmt_293_to_assign_stmt_792/slice_392_Update/ca
      -- 
    ca_948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_392_inst_ack_1, ack => maxPool4_CP_563_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	21 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	116 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 call_stmt_293_to_assign_stmt_792/slice_396_sample_start_
      -- CP-element group 114: 	 call_stmt_293_to_assign_stmt_792/slice_396_Sample/$entry
      -- CP-element group 114: 	 call_stmt_293_to_assign_stmt_792/slice_396_Sample/rr
      -- 
    rr_956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(114), ack => slice_396_inst_req_0); -- 
    maxPool4_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(21) & maxPool4_CP_563_elements(116);
      gj_maxPool4_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: marked-predecessors 
    -- CP-element group 115: 	117 
    -- CP-element group 115: 	164 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 call_stmt_293_to_assign_stmt_792/slice_396_update_start_
      -- CP-element group 115: 	 call_stmt_293_to_assign_stmt_792/slice_396_Update/$entry
      -- CP-element group 115: 	 call_stmt_293_to_assign_stmt_792/slice_396_Update/cr
      -- 
    cr_961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(115), ack => slice_396_inst_req_1); -- 
    maxPool4_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(117) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: marked-successors 
    -- CP-element group 116: 	19 
    -- CP-element group 116: 	114 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 call_stmt_293_to_assign_stmt_792/slice_396_sample_completed_
      -- CP-element group 116: 	 call_stmt_293_to_assign_stmt_792/slice_396_Sample/$exit
      -- CP-element group 116: 	 call_stmt_293_to_assign_stmt_792/slice_396_Sample/ra
      -- 
    ra_957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_396_inst_ack_0, ack => maxPool4_CP_563_elements(116)); -- 
    -- CP-element group 117:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	162 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	115 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 call_stmt_293_to_assign_stmt_792/slice_396_update_completed_
      -- CP-element group 117: 	 call_stmt_293_to_assign_stmt_792/slice_396_Update/$exit
      -- CP-element group 117: 	 call_stmt_293_to_assign_stmt_792/slice_396_Update/ca
      -- 
    ca_962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_396_inst_ack_1, ack => maxPool4_CP_563_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	21 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	120 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 call_stmt_293_to_assign_stmt_792/slice_400_sample_start_
      -- CP-element group 118: 	 call_stmt_293_to_assign_stmt_792/slice_400_Sample/$entry
      -- CP-element group 118: 	 call_stmt_293_to_assign_stmt_792/slice_400_Sample/rr
      -- 
    rr_970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(118), ack => slice_400_inst_req_0); -- 
    maxPool4_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(21) & maxPool4_CP_563_elements(120);
      gj_maxPool4_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	121 
    -- CP-element group 119: 	164 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 call_stmt_293_to_assign_stmt_792/slice_400_update_start_
      -- CP-element group 119: 	 call_stmt_293_to_assign_stmt_792/slice_400_Update/$entry
      -- CP-element group 119: 	 call_stmt_293_to_assign_stmt_792/slice_400_Update/cr
      -- 
    cr_975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(119), ack => slice_400_inst_req_1); -- 
    maxPool4_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(121) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: marked-successors 
    -- CP-element group 120: 	19 
    -- CP-element group 120: 	118 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 call_stmt_293_to_assign_stmt_792/slice_400_sample_completed_
      -- CP-element group 120: 	 call_stmt_293_to_assign_stmt_792/slice_400_Sample/$exit
      -- CP-element group 120: 	 call_stmt_293_to_assign_stmt_792/slice_400_Sample/ra
      -- 
    ra_971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_400_inst_ack_0, ack => maxPool4_CP_563_elements(120)); -- 
    -- CP-element group 121:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	162 
    -- CP-element group 121: marked-successors 
    -- CP-element group 121: 	119 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 call_stmt_293_to_assign_stmt_792/slice_400_update_completed_
      -- CP-element group 121: 	 call_stmt_293_to_assign_stmt_792/slice_400_Update/$exit
      -- CP-element group 121: 	 call_stmt_293_to_assign_stmt_792/slice_400_Update/ca
      -- 
    ca_976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_400_inst_ack_1, ack => maxPool4_CP_563_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	25 
    -- CP-element group 122: marked-predecessors 
    -- CP-element group 122: 	124 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 call_stmt_293_to_assign_stmt_792/slice_404_sample_start_
      -- CP-element group 122: 	 call_stmt_293_to_assign_stmt_792/slice_404_Sample/$entry
      -- CP-element group 122: 	 call_stmt_293_to_assign_stmt_792/slice_404_Sample/rr
      -- 
    rr_984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(122), ack => slice_404_inst_req_0); -- 
    maxPool4_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(25) & maxPool4_CP_563_elements(124);
      gj_maxPool4_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	164 
    -- CP-element group 123: 	168 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 call_stmt_293_to_assign_stmt_792/slice_404_update_start_
      -- CP-element group 123: 	 call_stmt_293_to_assign_stmt_792/slice_404_Update/$entry
      -- CP-element group 123: 	 call_stmt_293_to_assign_stmt_792/slice_404_Update/cr
      -- 
    cr_989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(123), ack => slice_404_inst_req_1); -- 
    maxPool4_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(125) & maxPool4_CP_563_elements(164) & maxPool4_CP_563_elements(168);
      gj_maxPool4_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: marked-successors 
    -- CP-element group 124: 	23 
    -- CP-element group 124: 	122 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 call_stmt_293_to_assign_stmt_792/slice_404_sample_completed_
      -- CP-element group 124: 	 call_stmt_293_to_assign_stmt_792/slice_404_Sample/$exit
      -- CP-element group 124: 	 call_stmt_293_to_assign_stmt_792/slice_404_Sample/ra
      -- 
    ra_985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_404_inst_ack_0, ack => maxPool4_CP_563_elements(124)); -- 
    -- CP-element group 125:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	162 
    -- CP-element group 125: 	166 
    -- CP-element group 125: marked-successors 
    -- CP-element group 125: 	123 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 call_stmt_293_to_assign_stmt_792/slice_404_update_completed_
      -- CP-element group 125: 	 call_stmt_293_to_assign_stmt_792/slice_404_Update/$exit
      -- CP-element group 125: 	 call_stmt_293_to_assign_stmt_792/slice_404_Update/ca
      -- 
    ca_990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_404_inst_ack_1, ack => maxPool4_CP_563_elements(125)); -- 
    -- CP-element group 126:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	25 
    -- CP-element group 126: marked-predecessors 
    -- CP-element group 126: 	128 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 call_stmt_293_to_assign_stmt_792/slice_408_sample_start_
      -- CP-element group 126: 	 call_stmt_293_to_assign_stmt_792/slice_408_Sample/$entry
      -- CP-element group 126: 	 call_stmt_293_to_assign_stmt_792/slice_408_Sample/rr
      -- 
    rr_998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(126), ack => slice_408_inst_req_0); -- 
    maxPool4_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(25) & maxPool4_CP_563_elements(128);
      gj_maxPool4_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: marked-predecessors 
    -- CP-element group 127: 	129 
    -- CP-element group 127: 	164 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 call_stmt_293_to_assign_stmt_792/slice_408_update_start_
      -- CP-element group 127: 	 call_stmt_293_to_assign_stmt_792/slice_408_Update/$entry
      -- CP-element group 127: 	 call_stmt_293_to_assign_stmt_792/slice_408_Update/cr
      -- 
    cr_1003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(127), ack => slice_408_inst_req_1); -- 
    maxPool4_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(129) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: marked-successors 
    -- CP-element group 128: 	23 
    -- CP-element group 128: 	126 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 call_stmt_293_to_assign_stmt_792/slice_408_sample_completed_
      -- CP-element group 128: 	 call_stmt_293_to_assign_stmt_792/slice_408_Sample/$exit
      -- CP-element group 128: 	 call_stmt_293_to_assign_stmt_792/slice_408_Sample/ra
      -- 
    ra_999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_408_inst_ack_0, ack => maxPool4_CP_563_elements(128)); -- 
    -- CP-element group 129:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	162 
    -- CP-element group 129: marked-successors 
    -- CP-element group 129: 	127 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 call_stmt_293_to_assign_stmt_792/slice_408_update_completed_
      -- CP-element group 129: 	 call_stmt_293_to_assign_stmt_792/slice_408_Update/$exit
      -- CP-element group 129: 	 call_stmt_293_to_assign_stmt_792/slice_408_Update/ca
      -- 
    ca_1004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_408_inst_ack_1, ack => maxPool4_CP_563_elements(129)); -- 
    -- CP-element group 130:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	25 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	132 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 call_stmt_293_to_assign_stmt_792/slice_412_sample_start_
      -- CP-element group 130: 	 call_stmt_293_to_assign_stmt_792/slice_412_Sample/$entry
      -- CP-element group 130: 	 call_stmt_293_to_assign_stmt_792/slice_412_Sample/rr
      -- 
    rr_1012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(130), ack => slice_412_inst_req_0); -- 
    maxPool4_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(25) & maxPool4_CP_563_elements(132);
      gj_maxPool4_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	133 
    -- CP-element group 131: 	164 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 call_stmt_293_to_assign_stmt_792/slice_412_update_start_
      -- CP-element group 131: 	 call_stmt_293_to_assign_stmt_792/slice_412_Update/$entry
      -- CP-element group 131: 	 call_stmt_293_to_assign_stmt_792/slice_412_Update/cr
      -- 
    cr_1017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(131), ack => slice_412_inst_req_1); -- 
    maxPool4_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(133) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: marked-successors 
    -- CP-element group 132: 	23 
    -- CP-element group 132: 	130 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 call_stmt_293_to_assign_stmt_792/slice_412_sample_completed_
      -- CP-element group 132: 	 call_stmt_293_to_assign_stmt_792/slice_412_Sample/$exit
      -- CP-element group 132: 	 call_stmt_293_to_assign_stmt_792/slice_412_Sample/ra
      -- 
    ra_1013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_412_inst_ack_0, ack => maxPool4_CP_563_elements(132)); -- 
    -- CP-element group 133:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	162 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	131 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 call_stmt_293_to_assign_stmt_792/slice_412_update_completed_
      -- CP-element group 133: 	 call_stmt_293_to_assign_stmt_792/slice_412_Update/$exit
      -- CP-element group 133: 	 call_stmt_293_to_assign_stmt_792/slice_412_Update/ca
      -- 
    ca_1018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_412_inst_ack_1, ack => maxPool4_CP_563_elements(133)); -- 
    -- CP-element group 134:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	25 
    -- CP-element group 134: marked-predecessors 
    -- CP-element group 134: 	136 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 call_stmt_293_to_assign_stmt_792/slice_416_sample_start_
      -- CP-element group 134: 	 call_stmt_293_to_assign_stmt_792/slice_416_Sample/$entry
      -- CP-element group 134: 	 call_stmt_293_to_assign_stmt_792/slice_416_Sample/rr
      -- 
    rr_1026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(134), ack => slice_416_inst_req_0); -- 
    maxPool4_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(25) & maxPool4_CP_563_elements(136);
      gj_maxPool4_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 135:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	137 
    -- CP-element group 135: 	164 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 call_stmt_293_to_assign_stmt_792/slice_416_update_start_
      -- CP-element group 135: 	 call_stmt_293_to_assign_stmt_792/slice_416_Update/$entry
      -- CP-element group 135: 	 call_stmt_293_to_assign_stmt_792/slice_416_Update/cr
      -- 
    cr_1031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(135), ack => slice_416_inst_req_1); -- 
    maxPool4_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(137) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: marked-successors 
    -- CP-element group 136: 	23 
    -- CP-element group 136: 	134 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 call_stmt_293_to_assign_stmt_792/slice_416_sample_completed_
      -- CP-element group 136: 	 call_stmt_293_to_assign_stmt_792/slice_416_Sample/$exit
      -- CP-element group 136: 	 call_stmt_293_to_assign_stmt_792/slice_416_Sample/ra
      -- 
    ra_1027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_416_inst_ack_0, ack => maxPool4_CP_563_elements(136)); -- 
    -- CP-element group 137:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	162 
    -- CP-element group 137: marked-successors 
    -- CP-element group 137: 	135 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 call_stmt_293_to_assign_stmt_792/slice_416_update_completed_
      -- CP-element group 137: 	 call_stmt_293_to_assign_stmt_792/slice_416_Update/$exit
      -- CP-element group 137: 	 call_stmt_293_to_assign_stmt_792/slice_416_Update/ca
      -- 
    ca_1032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_416_inst_ack_1, ack => maxPool4_CP_563_elements(137)); -- 
    -- CP-element group 138:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	25 
    -- CP-element group 138: marked-predecessors 
    -- CP-element group 138: 	140 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 call_stmt_293_to_assign_stmt_792/slice_420_sample_start_
      -- CP-element group 138: 	 call_stmt_293_to_assign_stmt_792/slice_420_Sample/$entry
      -- CP-element group 138: 	 call_stmt_293_to_assign_stmt_792/slice_420_Sample/rr
      -- 
    rr_1040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(138), ack => slice_420_inst_req_0); -- 
    maxPool4_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(25) & maxPool4_CP_563_elements(140);
      gj_maxPool4_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	141 
    -- CP-element group 139: 	164 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	141 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 call_stmt_293_to_assign_stmt_792/slice_420_update_start_
      -- CP-element group 139: 	 call_stmt_293_to_assign_stmt_792/slice_420_Update/$entry
      -- CP-element group 139: 	 call_stmt_293_to_assign_stmt_792/slice_420_Update/cr
      -- 
    cr_1045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(139), ack => slice_420_inst_req_1); -- 
    maxPool4_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(141) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140: marked-successors 
    -- CP-element group 140: 	23 
    -- CP-element group 140: 	138 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 call_stmt_293_to_assign_stmt_792/slice_420_sample_completed_
      -- CP-element group 140: 	 call_stmt_293_to_assign_stmt_792/slice_420_Sample/$exit
      -- CP-element group 140: 	 call_stmt_293_to_assign_stmt_792/slice_420_Sample/ra
      -- 
    ra_1041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_420_inst_ack_0, ack => maxPool4_CP_563_elements(140)); -- 
    -- CP-element group 141:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	162 
    -- CP-element group 141: marked-successors 
    -- CP-element group 141: 	139 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 call_stmt_293_to_assign_stmt_792/slice_420_update_completed_
      -- CP-element group 141: 	 call_stmt_293_to_assign_stmt_792/slice_420_Update/$exit
      -- CP-element group 141: 	 call_stmt_293_to_assign_stmt_792/slice_420_Update/ca
      -- 
    ca_1046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_420_inst_ack_1, ack => maxPool4_CP_563_elements(141)); -- 
    -- CP-element group 142:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	25 
    -- CP-element group 142: marked-predecessors 
    -- CP-element group 142: 	144 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 call_stmt_293_to_assign_stmt_792/slice_424_sample_start_
      -- CP-element group 142: 	 call_stmt_293_to_assign_stmt_792/slice_424_Sample/$entry
      -- CP-element group 142: 	 call_stmt_293_to_assign_stmt_792/slice_424_Sample/rr
      -- 
    rr_1054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(142), ack => slice_424_inst_req_0); -- 
    maxPool4_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(25) & maxPool4_CP_563_elements(144);
      gj_maxPool4_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	145 
    -- CP-element group 143: 	164 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 call_stmt_293_to_assign_stmt_792/slice_424_update_start_
      -- CP-element group 143: 	 call_stmt_293_to_assign_stmt_792/slice_424_Update/$entry
      -- CP-element group 143: 	 call_stmt_293_to_assign_stmt_792/slice_424_Update/cr
      -- 
    cr_1059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(143), ack => slice_424_inst_req_1); -- 
    maxPool4_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(145) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144: marked-successors 
    -- CP-element group 144: 	23 
    -- CP-element group 144: 	142 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 call_stmt_293_to_assign_stmt_792/slice_424_sample_completed_
      -- CP-element group 144: 	 call_stmt_293_to_assign_stmt_792/slice_424_Sample/$exit
      -- CP-element group 144: 	 call_stmt_293_to_assign_stmt_792/slice_424_Sample/ra
      -- 
    ra_1055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_424_inst_ack_0, ack => maxPool4_CP_563_elements(144)); -- 
    -- CP-element group 145:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	162 
    -- CP-element group 145: marked-successors 
    -- CP-element group 145: 	143 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 call_stmt_293_to_assign_stmt_792/slice_424_update_completed_
      -- CP-element group 145: 	 call_stmt_293_to_assign_stmt_792/slice_424_Update/$exit
      -- CP-element group 145: 	 call_stmt_293_to_assign_stmt_792/slice_424_Update/ca
      -- 
    ca_1060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_424_inst_ack_1, ack => maxPool4_CP_563_elements(145)); -- 
    -- CP-element group 146:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	25 
    -- CP-element group 146: marked-predecessors 
    -- CP-element group 146: 	148 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 call_stmt_293_to_assign_stmt_792/slice_428_sample_start_
      -- CP-element group 146: 	 call_stmt_293_to_assign_stmt_792/slice_428_Sample/$entry
      -- CP-element group 146: 	 call_stmt_293_to_assign_stmt_792/slice_428_Sample/rr
      -- 
    rr_1068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(146), ack => slice_428_inst_req_0); -- 
    maxPool4_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(25) & maxPool4_CP_563_elements(148);
      gj_maxPool4_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	149 
    -- CP-element group 147: 	164 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 call_stmt_293_to_assign_stmt_792/slice_428_update_start_
      -- CP-element group 147: 	 call_stmt_293_to_assign_stmt_792/slice_428_Update/$entry
      -- CP-element group 147: 	 call_stmt_293_to_assign_stmt_792/slice_428_Update/cr
      -- 
    cr_1073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(147), ack => slice_428_inst_req_1); -- 
    maxPool4_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(149) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148: marked-successors 
    -- CP-element group 148: 	23 
    -- CP-element group 148: 	146 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 call_stmt_293_to_assign_stmt_792/slice_428_sample_completed_
      -- CP-element group 148: 	 call_stmt_293_to_assign_stmt_792/slice_428_Sample/$exit
      -- CP-element group 148: 	 call_stmt_293_to_assign_stmt_792/slice_428_Sample/ra
      -- 
    ra_1069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_428_inst_ack_0, ack => maxPool4_CP_563_elements(148)); -- 
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	162 
    -- CP-element group 149: marked-successors 
    -- CP-element group 149: 	147 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 call_stmt_293_to_assign_stmt_792/slice_428_update_completed_
      -- CP-element group 149: 	 call_stmt_293_to_assign_stmt_792/slice_428_Update/$exit
      -- CP-element group 149: 	 call_stmt_293_to_assign_stmt_792/slice_428_Update/ca
      -- 
    ca_1074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_428_inst_ack_1, ack => maxPool4_CP_563_elements(149)); -- 
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	25 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	152 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 call_stmt_293_to_assign_stmt_792/slice_432_sample_start_
      -- CP-element group 150: 	 call_stmt_293_to_assign_stmt_792/slice_432_Sample/$entry
      -- CP-element group 150: 	 call_stmt_293_to_assign_stmt_792/slice_432_Sample/rr
      -- 
    rr_1082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(150), ack => slice_432_inst_req_0); -- 
    maxPool4_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(25) & maxPool4_CP_563_elements(152);
      gj_maxPool4_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	153 
    -- CP-element group 151: 	164 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 call_stmt_293_to_assign_stmt_792/slice_432_update_start_
      -- CP-element group 151: 	 call_stmt_293_to_assign_stmt_792/slice_432_Update/$entry
      -- CP-element group 151: 	 call_stmt_293_to_assign_stmt_792/slice_432_Update/cr
      -- 
    cr_1087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(151), ack => slice_432_inst_req_1); -- 
    maxPool4_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(153) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: marked-successors 
    -- CP-element group 152: 	23 
    -- CP-element group 152: 	150 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 call_stmt_293_to_assign_stmt_792/slice_432_sample_completed_
      -- CP-element group 152: 	 call_stmt_293_to_assign_stmt_792/slice_432_Sample/$exit
      -- CP-element group 152: 	 call_stmt_293_to_assign_stmt_792/slice_432_Sample/ra
      -- 
    ra_1083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_432_inst_ack_0, ack => maxPool4_CP_563_elements(152)); -- 
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	162 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	151 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 call_stmt_293_to_assign_stmt_792/slice_432_update_completed_
      -- CP-element group 153: 	 call_stmt_293_to_assign_stmt_792/slice_432_Update/$exit
      -- CP-element group 153: 	 call_stmt_293_to_assign_stmt_792/slice_432_Update/ca
      -- 
    ca_1088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_432_inst_ack_1, ack => maxPool4_CP_563_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	1 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_757_sample_start_
      -- CP-element group 154: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_757_Sample/$entry
      -- CP-element group 154: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_757_Sample/req
      -- 
    req_1096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(154), ack => W_index2_755_delayed_7_0_755_inst_req_0); -- 
    maxPool4_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(1) & maxPool4_CP_563_elements(156);
      gj_maxPool4_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	157 
    -- CP-element group 155: 	164 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_757_update_start_
      -- CP-element group 155: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_757_Update/$entry
      -- CP-element group 155: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_757_Update/req
      -- 
    req_1101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(155), ack => W_index2_755_delayed_7_0_755_inst_req_1); -- 
    maxPool4_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(157) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	8 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_757_sample_completed_
      -- CP-element group 156: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_757_Sample/$exit
      -- CP-element group 156: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_757_Sample/ack
      -- 
    ack_1097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index2_755_delayed_7_0_755_inst_ack_0, ack => maxPool4_CP_563_elements(156)); -- 
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	162 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	155 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_757_update_completed_
      -- CP-element group 157: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_757_Update/$exit
      -- CP-element group 157: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_757_Update/ack
      -- 
    ack_1102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index2_755_delayed_7_0_755_inst_ack_1, ack => maxPool4_CP_563_elements(157)); -- 
    -- CP-element group 158:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	1 
    -- CP-element group 158: marked-predecessors 
    -- CP-element group 158: 	160 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_760_sample_start_
      -- CP-element group 158: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_760_Sample/$entry
      -- CP-element group 158: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_760_Sample/req
      -- 
    req_1110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(158), ack => W_addr_756_delayed_7_0_758_inst_req_0); -- 
    maxPool4_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(1) & maxPool4_CP_563_elements(160);
      gj_maxPool4_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	161 
    -- CP-element group 159: 	164 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_760_update_start_
      -- CP-element group 159: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_760_Update/$entry
      -- CP-element group 159: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_760_Update/req
      -- 
    req_1115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(159), ack => W_addr_756_delayed_7_0_758_inst_req_1); -- 
    maxPool4_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(161) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160: marked-successors 
    -- CP-element group 160: 	2 
    -- CP-element group 160: 	158 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_760_sample_completed_
      -- CP-element group 160: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_760_Sample/$exit
      -- CP-element group 160: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_760_Sample/ack
      -- 
    ack_1111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_addr_756_delayed_7_0_758_inst_ack_0, ack => maxPool4_CP_563_elements(160)); -- 
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	159 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_760_update_completed_
      -- CP-element group 161: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_760_Update/$exit
      -- CP-element group 161: 	 call_stmt_293_to_assign_stmt_792/assign_stmt_760_Update/ack
      -- 
    ack_1116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_addr_756_delayed_7_0_758_inst_ack_1, ack => maxPool4_CP_563_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	41 
    -- CP-element group 162: 	45 
    -- CP-element group 162: 	49 
    -- CP-element group 162: 	53 
    -- CP-element group 162: 	57 
    -- CP-element group 162: 	61 
    -- CP-element group 162: 	65 
    -- CP-element group 162: 	69 
    -- CP-element group 162: 	73 
    -- CP-element group 162: 	77 
    -- CP-element group 162: 	81 
    -- CP-element group 162: 	37 
    -- CP-element group 162: 	29 
    -- CP-element group 162: 	33 
    -- CP-element group 162: 	85 
    -- CP-element group 162: 	89 
    -- CP-element group 162: 	93 
    -- CP-element group 162: 	97 
    -- CP-element group 162: 	101 
    -- CP-element group 162: 	105 
    -- CP-element group 162: 	109 
    -- CP-element group 162: 	113 
    -- CP-element group 162: 	117 
    -- CP-element group 162: 	121 
    -- CP-element group 162: 	125 
    -- CP-element group 162: 	129 
    -- CP-element group 162: 	133 
    -- CP-element group 162: 	137 
    -- CP-element group 162: 	141 
    -- CP-element group 162: 	145 
    -- CP-element group 162: 	149 
    -- CP-element group 162: 	153 
    -- CP-element group 162: 	157 
    -- CP-element group 162: 	161 
    -- CP-element group 162: marked-predecessors 
    -- CP-element group 162: 	164 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	164 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 call_stmt_293_to_assign_stmt_792/call_stmt_788_sample_start_
      -- CP-element group 162: 	 call_stmt_293_to_assign_stmt_792/call_stmt_788_Sample/$entry
      -- CP-element group 162: 	 call_stmt_293_to_assign_stmt_792/call_stmt_788_Sample/crr
      -- 
    crr_1124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(162), ack => call_stmt_788_call_req_0); -- 
    maxPool4_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 34) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1,28 => 1,29 => 1,30 => 1,31 => 1,32 => 1,33 => 1,34 => 1);
      constant place_markings: IntegerArray(0 to 34)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0,26 => 0,27 => 0,28 => 0,29 => 0,30 => 0,31 => 0,32 => 0,33 => 0,34 => 1);
      constant place_delays: IntegerArray(0 to 34) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0,26 => 0,27 => 0,28 => 0,29 => 0,30 => 0,31 => 0,32 => 0,33 => 0,34 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 35); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(41) & maxPool4_CP_563_elements(45) & maxPool4_CP_563_elements(49) & maxPool4_CP_563_elements(53) & maxPool4_CP_563_elements(57) & maxPool4_CP_563_elements(61) & maxPool4_CP_563_elements(65) & maxPool4_CP_563_elements(69) & maxPool4_CP_563_elements(73) & maxPool4_CP_563_elements(77) & maxPool4_CP_563_elements(81) & maxPool4_CP_563_elements(37) & maxPool4_CP_563_elements(29) & maxPool4_CP_563_elements(33) & maxPool4_CP_563_elements(85) & maxPool4_CP_563_elements(89) & maxPool4_CP_563_elements(93) & maxPool4_CP_563_elements(97) & maxPool4_CP_563_elements(101) & maxPool4_CP_563_elements(105) & maxPool4_CP_563_elements(109) & maxPool4_CP_563_elements(113) & maxPool4_CP_563_elements(117) & maxPool4_CP_563_elements(121) & maxPool4_CP_563_elements(125) & maxPool4_CP_563_elements(129) & maxPool4_CP_563_elements(133) & maxPool4_CP_563_elements(137) & maxPool4_CP_563_elements(141) & maxPool4_CP_563_elements(145) & maxPool4_CP_563_elements(149) & maxPool4_CP_563_elements(153) & maxPool4_CP_563_elements(157) & maxPool4_CP_563_elements(161) & maxPool4_CP_563_elements(164);
      gj_maxPool4_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 35, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 call_stmt_293_to_assign_stmt_792/call_stmt_788_update_start_
      -- CP-element group 163: 	 call_stmt_293_to_assign_stmt_792/call_stmt_788_Update/$entry
      -- CP-element group 163: 	 call_stmt_293_to_assign_stmt_792/call_stmt_788_Update/ccr
      -- 
    ccr_1129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(163), ack => call_stmt_788_call_req_1); -- 
    maxPool4_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_563_elements(165);
      gj_maxPool4_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164: marked-successors 
    -- CP-element group 164: 	39 
    -- CP-element group 164: 	43 
    -- CP-element group 164: 	47 
    -- CP-element group 164: 	51 
    -- CP-element group 164: 	55 
    -- CP-element group 164: 	59 
    -- CP-element group 164: 	63 
    -- CP-element group 164: 	67 
    -- CP-element group 164: 	71 
    -- CP-element group 164: 	75 
    -- CP-element group 164: 	79 
    -- CP-element group 164: 	83 
    -- CP-element group 164: 	35 
    -- CP-element group 164: 	27 
    -- CP-element group 164: 	31 
    -- CP-element group 164: 	87 
    -- CP-element group 164: 	91 
    -- CP-element group 164: 	95 
    -- CP-element group 164: 	99 
    -- CP-element group 164: 	103 
    -- CP-element group 164: 	107 
    -- CP-element group 164: 	111 
    -- CP-element group 164: 	115 
    -- CP-element group 164: 	119 
    -- CP-element group 164: 	123 
    -- CP-element group 164: 	127 
    -- CP-element group 164: 	131 
    -- CP-element group 164: 	135 
    -- CP-element group 164: 	139 
    -- CP-element group 164: 	143 
    -- CP-element group 164: 	147 
    -- CP-element group 164: 	151 
    -- CP-element group 164: 	155 
    -- CP-element group 164: 	159 
    -- CP-element group 164: 	162 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 call_stmt_293_to_assign_stmt_792/call_stmt_788_sample_completed_
      -- CP-element group 164: 	 call_stmt_293_to_assign_stmt_792/call_stmt_788_Sample/$exit
      -- CP-element group 164: 	 call_stmt_293_to_assign_stmt_792/call_stmt_788_Sample/cra
      -- 
    cra_1125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_788_call_ack_0, ack => maxPool4_CP_563_elements(164)); -- 
    -- CP-element group 165:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	170 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	163 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 call_stmt_293_to_assign_stmt_792/call_stmt_788_update_completed_
      -- CP-element group 165: 	 call_stmt_293_to_assign_stmt_792/call_stmt_788_Update/$exit
      -- CP-element group 165: 	 call_stmt_293_to_assign_stmt_792/call_stmt_788_Update/cca
      -- 
    cca_1130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_788_call_ack_1, ack => maxPool4_CP_563_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	61 
    -- CP-element group 166: 	29 
    -- CP-element group 166: 	93 
    -- CP-element group 166: 	125 
    -- CP-element group 166: marked-predecessors 
    -- CP-element group 166: 	168 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	168 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 call_stmt_293_to_assign_stmt_792/type_cast_791_sample_start_
      -- CP-element group 166: 	 call_stmt_293_to_assign_stmt_792/type_cast_791_Sample/$entry
      -- CP-element group 166: 	 call_stmt_293_to_assign_stmt_792/type_cast_791_Sample/rr
      -- 
    rr_1138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(166), ack => type_cast_791_inst_req_0); -- 
    maxPool4_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(61) & maxPool4_CP_563_elements(29) & maxPool4_CP_563_elements(93) & maxPool4_CP_563_elements(125) & maxPool4_CP_563_elements(168);
      gj_maxPool4_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	9 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	169 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 call_stmt_293_to_assign_stmt_792/type_cast_791_update_start_
      -- CP-element group 167: 	 call_stmt_293_to_assign_stmt_792/type_cast_791_Update/$entry
      -- CP-element group 167: 	 call_stmt_293_to_assign_stmt_792/type_cast_791_Update/cr
      -- 
    cr_1143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_563_elements(167), ack => type_cast_791_inst_req_1); -- 
    maxPool4_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(9) & maxPool4_CP_563_elements(169);
      gj_maxPool4_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168: marked-successors 
    -- CP-element group 168: 	59 
    -- CP-element group 168: 	27 
    -- CP-element group 168: 	91 
    -- CP-element group 168: 	123 
    -- CP-element group 168: 	166 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 call_stmt_293_to_assign_stmt_792/type_cast_791_sample_completed_
      -- CP-element group 168: 	 call_stmt_293_to_assign_stmt_792/type_cast_791_Sample/$exit
      -- CP-element group 168: 	 call_stmt_293_to_assign_stmt_792/type_cast_791_Sample/ra
      -- 
    ra_1139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_791_inst_ack_0, ack => maxPool4_CP_563_elements(168)); -- 
    -- CP-element group 169:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169: marked-successors 
    -- CP-element group 169: 	167 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 call_stmt_293_to_assign_stmt_792/type_cast_791_update_completed_
      -- CP-element group 169: 	 call_stmt_293_to_assign_stmt_792/type_cast_791_Update/$exit
      -- CP-element group 169: 	 call_stmt_293_to_assign_stmt_792/type_cast_791_Update/ca
      -- 
    ca_1144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_791_inst_ack_1, ack => maxPool4_CP_563_elements(169)); -- 
    -- CP-element group 170:  join  transition  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	165 
    -- CP-element group 170: 	169 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	179 
    -- CP-element group 170:  members (1) 
      -- CP-element group 170: 	 call_stmt_293_to_assign_stmt_792/$exit
      -- 
    maxPool4_cp_element_group_170: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_170"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_563_elements(165) & maxPool4_CP_563_elements(169);
      gj_maxPool4_cp_element_group_170 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_563_elements(170), clk => clk, reset => reset); --
    end block;
    -- CP-element group 171:  place  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	2 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (1) 
      -- CP-element group 171: 	 addr_update_enable
      -- 
    maxPool4_CP_563_elements(171) <= maxPool4_CP_563_elements(2);
    -- CP-element group 172:  place  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	3 
    -- CP-element group 172: successors 
    -- CP-element group 172:  members (1) 
      -- CP-element group 172: 	 addr1_update_enable
      -- 
    maxPool4_CP_563_elements(172) <= maxPool4_CP_563_elements(3);
    -- CP-element group 173:  place  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	4 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (1) 
      -- CP-element group 173: 	 addr2_update_enable
      -- 
    maxPool4_CP_563_elements(173) <= maxPool4_CP_563_elements(4);
    -- CP-element group 174:  place  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	5 
    -- CP-element group 174: successors 
    -- CP-element group 174:  members (1) 
      -- CP-element group 174: 	 addr3_update_enable
      -- 
    maxPool4_CP_563_elements(174) <= maxPool4_CP_563_elements(5);
    -- CP-element group 175:  place  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	6 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (1) 
      -- CP-element group 175: 	 addr4_update_enable
      -- 
    maxPool4_CP_563_elements(175) <= maxPool4_CP_563_elements(6);
    -- CP-element group 176:  place  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	7 
    -- CP-element group 176: successors 
    -- CP-element group 176:  members (1) 
      -- CP-element group 176: 	 index1_update_enable
      -- 
    maxPool4_CP_563_elements(176) <= maxPool4_CP_563_elements(7);
    -- CP-element group 177:  place  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	8 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (1) 
      -- CP-element group 177: 	 index2_update_enable
      -- 
    maxPool4_CP_563_elements(177) <= maxPool4_CP_563_elements(8);
    -- CP-element group 178:  place  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	9 
    -- CP-element group 178:  members (1) 
      -- CP-element group 178: 	 output_update_enable
      -- 
    -- CP-element group 179:  transition  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	170 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (1) 
      -- CP-element group 179: 	 $exit
      -- 
    maxPool4_CP_563_elements(179) <= maxPool4_CP_563_elements(170);
    --  hookup: inputs to control-path 
    maxPool4_CP_563_elements(178) <= output_update_enable;
    -- hookup: output from control-path 
    addr_update_enable <= maxPool4_CP_563_elements(171);
    addr1_update_enable <= maxPool4_CP_563_elements(172);
    addr2_update_enable <= maxPool4_CP_563_elements(173);
    addr3_update_enable <= maxPool4_CP_563_elements(174);
    addr4_update_enable <= maxPool4_CP_563_elements(175);
    index1_update_enable <= maxPool4_CP_563_elements(176);
    index2_update_enable <= maxPool4_CP_563_elements(177);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u16_u32_774_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_785_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u32_u64_786_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u8_u16_767_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_773_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_779_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_784_wire : std_logic_vector(15 downto 0);
    signal SGT_i8_u1_566_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_574_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_582_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_590_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_598_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_606_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_614_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_622_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_630_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_638_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_646_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_654_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_662_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_670_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_678_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_686_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_694_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_702_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_710_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_718_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_726_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_734_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_742_wire : std_logic_vector(0 downto 0);
    signal SGT_i8_u1_750_wire : std_logic_vector(0 downto 0);
    signal a11_438 : std_logic_vector(7 downto 0);
    signal a12_442 : std_logic_vector(7 downto 0);
    signal a13_446 : std_logic_vector(7 downto 0);
    signal a14_450 : std_logic_vector(7 downto 0);
    signal a15_454 : std_logic_vector(7 downto 0);
    signal a16_458 : std_logic_vector(7 downto 0);
    signal a17_462 : std_logic_vector(7 downto 0);
    signal a18_466 : std_logic_vector(7 downto 0);
    signal a21_470 : std_logic_vector(7 downto 0);
    signal a22_474 : std_logic_vector(7 downto 0);
    signal a23_478 : std_logic_vector(7 downto 0);
    signal a24_482 : std_logic_vector(7 downto 0);
    signal a25_486 : std_logic_vector(7 downto 0);
    signal a26_490 : std_logic_vector(7 downto 0);
    signal a27_494 : std_logic_vector(7 downto 0);
    signal a28_498 : std_logic_vector(7 downto 0);
    signal a31_502 : std_logic_vector(7 downto 0);
    signal a32_506 : std_logic_vector(7 downto 0);
    signal a33_510 : std_logic_vector(7 downto 0);
    signal a34_514 : std_logic_vector(7 downto 0);
    signal a35_518 : std_logic_vector(7 downto 0);
    signal a36_522 : std_logic_vector(7 downto 0);
    signal a37_526 : std_logic_vector(7 downto 0);
    signal a38_530 : std_logic_vector(7 downto 0);
    signal a41_534 : std_logic_vector(7 downto 0);
    signal a42_538 : std_logic_vector(7 downto 0);
    signal a43_542 : std_logic_vector(7 downto 0);
    signal a44_546 : std_logic_vector(7 downto 0);
    signal a45_550 : std_logic_vector(7 downto 0);
    signal a46_554 : std_logic_vector(7 downto 0);
    signal a47_558 : std_logic_vector(7 downto 0);
    signal a48_562 : std_logic_vector(7 downto 0);
    signal addr_756_delayed_7_0_760 : std_logic_vector(31 downto 0);
    signal c1_293 : std_logic_vector(63 downto 0);
    signal c2_297 : std_logic_vector(63 downto 0);
    signal c3_301 : std_logic_vector(63 downto 0);
    signal c4_305 : std_logic_vector(63 downto 0);
    signal d1_788 : std_logic_vector(0 downto 0);
    signal index2_755_delayed_7_0_757 : std_logic_vector(7 downto 0);
    signal out1_586 : std_logic_vector(7 downto 0);
    signal out2_610 : std_logic_vector(7 downto 0);
    signal out3_634 : std_logic_vector(7 downto 0);
    signal out4_658 : std_logic_vector(7 downto 0);
    signal out5_682 : std_logic_vector(7 downto 0);
    signal out6_706 : std_logic_vector(7 downto 0);
    signal out7_730 : std_logic_vector(7 downto 0);
    signal out8_754 : std_logic_vector(7 downto 0);
    signal sliced_v11_309 : std_logic_vector(7 downto 0);
    signal sliced_v12_313 : std_logic_vector(7 downto 0);
    signal sliced_v13_317 : std_logic_vector(7 downto 0);
    signal sliced_v14_321 : std_logic_vector(7 downto 0);
    signal sliced_v15_325 : std_logic_vector(7 downto 0);
    signal sliced_v16_329 : std_logic_vector(7 downto 0);
    signal sliced_v17_333 : std_logic_vector(7 downto 0);
    signal sliced_v18_337 : std_logic_vector(7 downto 0);
    signal sliced_v21_341 : std_logic_vector(7 downto 0);
    signal sliced_v22_345 : std_logic_vector(7 downto 0);
    signal sliced_v23_349 : std_logic_vector(7 downto 0);
    signal sliced_v24_353 : std_logic_vector(7 downto 0);
    signal sliced_v25_357 : std_logic_vector(7 downto 0);
    signal sliced_v26_361 : std_logic_vector(7 downto 0);
    signal sliced_v27_365 : std_logic_vector(7 downto 0);
    signal sliced_v28_369 : std_logic_vector(7 downto 0);
    signal sliced_v31_373 : std_logic_vector(7 downto 0);
    signal sliced_v32_377 : std_logic_vector(7 downto 0);
    signal sliced_v33_381 : std_logic_vector(7 downto 0);
    signal sliced_v34_385 : std_logic_vector(7 downto 0);
    signal sliced_v35_389 : std_logic_vector(7 downto 0);
    signal sliced_v36_393 : std_logic_vector(7 downto 0);
    signal sliced_v37_397 : std_logic_vector(7 downto 0);
    signal sliced_v38_401 : std_logic_vector(7 downto 0);
    signal sliced_v41_405 : std_logic_vector(7 downto 0);
    signal sliced_v42_409 : std_logic_vector(7 downto 0);
    signal sliced_v43_413 : std_logic_vector(7 downto 0);
    signal sliced_v44_417 : std_logic_vector(7 downto 0);
    signal sliced_v45_421 : std_logic_vector(7 downto 0);
    signal sliced_v46_425 : std_logic_vector(7 downto 0);
    signal sliced_v47_429 : std_logic_vector(7 downto 0);
    signal sliced_v48_433 : std_logic_vector(7 downto 0);
    signal t11_570 : std_logic_vector(7 downto 0);
    signal t12_578 : std_logic_vector(7 downto 0);
    signal t21_594 : std_logic_vector(7 downto 0);
    signal t22_602 : std_logic_vector(7 downto 0);
    signal t31_618 : std_logic_vector(7 downto 0);
    signal t32_626 : std_logic_vector(7 downto 0);
    signal t41_642 : std_logic_vector(7 downto 0);
    signal t42_650 : std_logic_vector(7 downto 0);
    signal t51_666 : std_logic_vector(7 downto 0);
    signal t52_674 : std_logic_vector(7 downto 0);
    signal t61_690 : std_logic_vector(7 downto 0);
    signal t62_698 : std_logic_vector(7 downto 0);
    signal t71_714 : std_logic_vector(7 downto 0);
    signal t72_722 : std_logic_vector(7 downto 0);
    signal t81_738 : std_logic_vector(7 downto 0);
    signal t82_746 : std_logic_vector(7 downto 0);
    signal type_cast_764_wire : std_logic_vector(7 downto 0);
    signal type_cast_766_wire : std_logic_vector(7 downto 0);
    signal type_cast_770_wire : std_logic_vector(7 downto 0);
    signal type_cast_772_wire : std_logic_vector(7 downto 0);
    signal type_cast_776_wire : std_logic_vector(7 downto 0);
    signal type_cast_778_wire : std_logic_vector(7 downto 0);
    signal type_cast_781_wire : std_logic_vector(7 downto 0);
    signal type_cast_783_wire : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    -- flow-through select operator MUX_569_inst
    t11_570 <= a11_438 when (SGT_i8_u1_566_wire(0) /=  '0') else a21_470;
    -- flow-through select operator MUX_577_inst
    t12_578 <= a31_502 when (SGT_i8_u1_574_wire(0) /=  '0') else a41_534;
    -- flow-through select operator MUX_585_inst
    out1_586 <= t11_570 when (SGT_i8_u1_582_wire(0) /=  '0') else t12_578;
    -- flow-through select operator MUX_593_inst
    t21_594 <= a12_442 when (SGT_i8_u1_590_wire(0) /=  '0') else a22_474;
    -- flow-through select operator MUX_601_inst
    t22_602 <= a32_506 when (SGT_i8_u1_598_wire(0) /=  '0') else a42_538;
    -- flow-through select operator MUX_609_inst
    out2_610 <= t21_594 when (SGT_i8_u1_606_wire(0) /=  '0') else t22_602;
    -- flow-through select operator MUX_617_inst
    t31_618 <= a13_446 when (SGT_i8_u1_614_wire(0) /=  '0') else a23_478;
    -- flow-through select operator MUX_625_inst
    t32_626 <= a33_510 when (SGT_i8_u1_622_wire(0) /=  '0') else a43_542;
    -- flow-through select operator MUX_633_inst
    out3_634 <= t31_618 when (SGT_i8_u1_630_wire(0) /=  '0') else t32_626;
    -- flow-through select operator MUX_641_inst
    t41_642 <= a14_450 when (SGT_i8_u1_638_wire(0) /=  '0') else a24_482;
    -- flow-through select operator MUX_649_inst
    t42_650 <= a34_514 when (SGT_i8_u1_646_wire(0) /=  '0') else a44_546;
    -- flow-through select operator MUX_657_inst
    out4_658 <= t41_642 when (SGT_i8_u1_654_wire(0) /=  '0') else t42_650;
    -- flow-through select operator MUX_665_inst
    t51_666 <= a15_454 when (SGT_i8_u1_662_wire(0) /=  '0') else a25_486;
    -- flow-through select operator MUX_673_inst
    t52_674 <= a35_518 when (SGT_i8_u1_670_wire(0) /=  '0') else a45_550;
    -- flow-through select operator MUX_681_inst
    out5_682 <= t51_666 when (SGT_i8_u1_678_wire(0) /=  '0') else t52_674;
    -- flow-through select operator MUX_689_inst
    t61_690 <= a16_458 when (SGT_i8_u1_686_wire(0) /=  '0') else a26_490;
    -- flow-through select operator MUX_697_inst
    t62_698 <= a36_522 when (SGT_i8_u1_694_wire(0) /=  '0') else a46_554;
    -- flow-through select operator MUX_705_inst
    out6_706 <= t61_690 when (SGT_i8_u1_702_wire(0) /=  '0') else t62_698;
    -- flow-through select operator MUX_713_inst
    t71_714 <= a17_462 when (SGT_i8_u1_710_wire(0) /=  '0') else a27_494;
    -- flow-through select operator MUX_721_inst
    t72_722 <= a37_526 when (SGT_i8_u1_718_wire(0) /=  '0') else a47_558;
    -- flow-through select operator MUX_729_inst
    out7_730 <= t71_714 when (SGT_i8_u1_726_wire(0) /=  '0') else t72_722;
    -- flow-through select operator MUX_737_inst
    t81_738 <= a18_466 when (SGT_i8_u1_734_wire(0) /=  '0') else a28_498;
    -- flow-through select operator MUX_745_inst
    t82_746 <= a38_530 when (SGT_i8_u1_742_wire(0) /=  '0') else a48_562;
    -- flow-through select operator MUX_753_inst
    out8_754 <= t81_738 when (SGT_i8_u1_750_wire(0) /=  '0') else t82_746;
    slice_308_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_308_inst_req_0;
      slice_308_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_308_inst_req_1;
      slice_308_inst_ack_1<= update_ack(0);
      slice_308_inst: SliceSplitProtocol generic map(name => "slice_308_inst", in_data_width => 64, high_index => 63, low_index => 56, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_293, dout => sliced_v11_309, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_312_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_312_inst_req_0;
      slice_312_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_312_inst_req_1;
      slice_312_inst_ack_1<= update_ack(0);
      slice_312_inst: SliceSplitProtocol generic map(name => "slice_312_inst", in_data_width => 64, high_index => 55, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_293, dout => sliced_v12_313, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_316_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_316_inst_req_0;
      slice_316_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_316_inst_req_1;
      slice_316_inst_ack_1<= update_ack(0);
      slice_316_inst: SliceSplitProtocol generic map(name => "slice_316_inst", in_data_width => 64, high_index => 47, low_index => 40, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_293, dout => sliced_v13_317, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_320_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_320_inst_req_0;
      slice_320_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_320_inst_req_1;
      slice_320_inst_ack_1<= update_ack(0);
      slice_320_inst: SliceSplitProtocol generic map(name => "slice_320_inst", in_data_width => 64, high_index => 39, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_293, dout => sliced_v14_321, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_324_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_324_inst_req_0;
      slice_324_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_324_inst_req_1;
      slice_324_inst_ack_1<= update_ack(0);
      slice_324_inst: SliceSplitProtocol generic map(name => "slice_324_inst", in_data_width => 64, high_index => 31, low_index => 24, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_293, dout => sliced_v15_325, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_328_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_328_inst_req_0;
      slice_328_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_328_inst_req_1;
      slice_328_inst_ack_1<= update_ack(0);
      slice_328_inst: SliceSplitProtocol generic map(name => "slice_328_inst", in_data_width => 64, high_index => 23, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_293, dout => sliced_v16_329, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_332_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_332_inst_req_0;
      slice_332_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_332_inst_req_1;
      slice_332_inst_ack_1<= update_ack(0);
      slice_332_inst: SliceSplitProtocol generic map(name => "slice_332_inst", in_data_width => 64, high_index => 15, low_index => 8, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_293, dout => sliced_v17_333, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_336_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_336_inst_req_0;
      slice_336_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_336_inst_req_1;
      slice_336_inst_ack_1<= update_ack(0);
      slice_336_inst: SliceSplitProtocol generic map(name => "slice_336_inst", in_data_width => 64, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_293, dout => sliced_v18_337, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_340_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_340_inst_req_0;
      slice_340_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_340_inst_req_1;
      slice_340_inst_ack_1<= update_ack(0);
      slice_340_inst: SliceSplitProtocol generic map(name => "slice_340_inst", in_data_width => 64, high_index => 63, low_index => 56, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_297, dout => sliced_v21_341, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_344_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_344_inst_req_0;
      slice_344_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_344_inst_req_1;
      slice_344_inst_ack_1<= update_ack(0);
      slice_344_inst: SliceSplitProtocol generic map(name => "slice_344_inst", in_data_width => 64, high_index => 55, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_297, dout => sliced_v22_345, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_348_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_348_inst_req_0;
      slice_348_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_348_inst_req_1;
      slice_348_inst_ack_1<= update_ack(0);
      slice_348_inst: SliceSplitProtocol generic map(name => "slice_348_inst", in_data_width => 64, high_index => 47, low_index => 40, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_297, dout => sliced_v23_349, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_352_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_352_inst_req_0;
      slice_352_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_352_inst_req_1;
      slice_352_inst_ack_1<= update_ack(0);
      slice_352_inst: SliceSplitProtocol generic map(name => "slice_352_inst", in_data_width => 64, high_index => 39, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_297, dout => sliced_v24_353, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_356_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_356_inst_req_0;
      slice_356_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_356_inst_req_1;
      slice_356_inst_ack_1<= update_ack(0);
      slice_356_inst: SliceSplitProtocol generic map(name => "slice_356_inst", in_data_width => 64, high_index => 31, low_index => 24, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_297, dout => sliced_v25_357, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_360_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_360_inst_req_0;
      slice_360_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_360_inst_req_1;
      slice_360_inst_ack_1<= update_ack(0);
      slice_360_inst: SliceSplitProtocol generic map(name => "slice_360_inst", in_data_width => 64, high_index => 23, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_297, dout => sliced_v26_361, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_364_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_364_inst_req_0;
      slice_364_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_364_inst_req_1;
      slice_364_inst_ack_1<= update_ack(0);
      slice_364_inst: SliceSplitProtocol generic map(name => "slice_364_inst", in_data_width => 64, high_index => 15, low_index => 8, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_297, dout => sliced_v27_365, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_368_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_368_inst_req_0;
      slice_368_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_368_inst_req_1;
      slice_368_inst_ack_1<= update_ack(0);
      slice_368_inst: SliceSplitProtocol generic map(name => "slice_368_inst", in_data_width => 64, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_297, dout => sliced_v28_369, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_372_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_372_inst_req_0;
      slice_372_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_372_inst_req_1;
      slice_372_inst_ack_1<= update_ack(0);
      slice_372_inst: SliceSplitProtocol generic map(name => "slice_372_inst", in_data_width => 64, high_index => 63, low_index => 56, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_301, dout => sliced_v31_373, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_376_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_376_inst_req_0;
      slice_376_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_376_inst_req_1;
      slice_376_inst_ack_1<= update_ack(0);
      slice_376_inst: SliceSplitProtocol generic map(name => "slice_376_inst", in_data_width => 64, high_index => 55, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_301, dout => sliced_v32_377, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_380_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_380_inst_req_0;
      slice_380_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_380_inst_req_1;
      slice_380_inst_ack_1<= update_ack(0);
      slice_380_inst: SliceSplitProtocol generic map(name => "slice_380_inst", in_data_width => 64, high_index => 47, low_index => 40, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_301, dout => sliced_v33_381, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_384_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_384_inst_req_0;
      slice_384_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_384_inst_req_1;
      slice_384_inst_ack_1<= update_ack(0);
      slice_384_inst: SliceSplitProtocol generic map(name => "slice_384_inst", in_data_width => 64, high_index => 39, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_301, dout => sliced_v34_385, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_388_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_388_inst_req_0;
      slice_388_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_388_inst_req_1;
      slice_388_inst_ack_1<= update_ack(0);
      slice_388_inst: SliceSplitProtocol generic map(name => "slice_388_inst", in_data_width => 64, high_index => 31, low_index => 24, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_301, dout => sliced_v35_389, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_392_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_392_inst_req_0;
      slice_392_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_392_inst_req_1;
      slice_392_inst_ack_1<= update_ack(0);
      slice_392_inst: SliceSplitProtocol generic map(name => "slice_392_inst", in_data_width => 64, high_index => 23, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_301, dout => sliced_v36_393, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_396_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_396_inst_req_0;
      slice_396_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_396_inst_req_1;
      slice_396_inst_ack_1<= update_ack(0);
      slice_396_inst: SliceSplitProtocol generic map(name => "slice_396_inst", in_data_width => 64, high_index => 15, low_index => 8, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_301, dout => sliced_v37_397, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_400_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_400_inst_req_0;
      slice_400_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_400_inst_req_1;
      slice_400_inst_ack_1<= update_ack(0);
      slice_400_inst: SliceSplitProtocol generic map(name => "slice_400_inst", in_data_width => 64, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_301, dout => sliced_v38_401, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_404_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_404_inst_req_0;
      slice_404_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_404_inst_req_1;
      slice_404_inst_ack_1<= update_ack(0);
      slice_404_inst: SliceSplitProtocol generic map(name => "slice_404_inst", in_data_width => 64, high_index => 63, low_index => 56, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_305, dout => sliced_v41_405, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_408_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_408_inst_req_0;
      slice_408_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_408_inst_req_1;
      slice_408_inst_ack_1<= update_ack(0);
      slice_408_inst: SliceSplitProtocol generic map(name => "slice_408_inst", in_data_width => 64, high_index => 55, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_305, dout => sliced_v42_409, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_412_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_412_inst_req_0;
      slice_412_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_412_inst_req_1;
      slice_412_inst_ack_1<= update_ack(0);
      slice_412_inst: SliceSplitProtocol generic map(name => "slice_412_inst", in_data_width => 64, high_index => 47, low_index => 40, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_305, dout => sliced_v43_413, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_416_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_416_inst_req_0;
      slice_416_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_416_inst_req_1;
      slice_416_inst_ack_1<= update_ack(0);
      slice_416_inst: SliceSplitProtocol generic map(name => "slice_416_inst", in_data_width => 64, high_index => 39, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_305, dout => sliced_v44_417, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_420_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_420_inst_req_0;
      slice_420_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_420_inst_req_1;
      slice_420_inst_ack_1<= update_ack(0);
      slice_420_inst: SliceSplitProtocol generic map(name => "slice_420_inst", in_data_width => 64, high_index => 31, low_index => 24, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_305, dout => sliced_v45_421, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_424_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_424_inst_req_0;
      slice_424_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_424_inst_req_1;
      slice_424_inst_ack_1<= update_ack(0);
      slice_424_inst: SliceSplitProtocol generic map(name => "slice_424_inst", in_data_width => 64, high_index => 23, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_305, dout => sliced_v46_425, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_428_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_428_inst_req_0;
      slice_428_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_428_inst_req_1;
      slice_428_inst_ack_1<= update_ack(0);
      slice_428_inst: SliceSplitProtocol generic map(name => "slice_428_inst", in_data_width => 64, high_index => 15, low_index => 8, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_305, dout => sliced_v47_429, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_432_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_432_inst_req_0;
      slice_432_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_432_inst_req_1;
      slice_432_inst_ack_1<= update_ack(0);
      slice_432_inst: SliceSplitProtocol generic map(name => "slice_432_inst", in_data_width => 64, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_305, dout => sliced_v48_433, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_addr_756_delayed_7_0_758_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_addr_756_delayed_7_0_758_inst_req_0;
      W_addr_756_delayed_7_0_758_inst_ack_0<= wack(0);
      rreq(0) <= W_addr_756_delayed_7_0_758_inst_req_1;
      W_addr_756_delayed_7_0_758_inst_ack_1<= rack(0);
      W_addr_756_delayed_7_0_758_inst : InterlockBuffer generic map ( -- 
        name => "W_addr_756_delayed_7_0_758_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => addr_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => addr_756_delayed_7_0_760,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_index2_755_delayed_7_0_755_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_index2_755_delayed_7_0_755_inst_req_0;
      W_index2_755_delayed_7_0_755_inst_ack_0<= wack(0);
      rreq(0) <= W_index2_755_delayed_7_0_755_inst_req_1;
      W_index2_755_delayed_7_0_755_inst_ack_1<= rack(0);
      W_index2_755_delayed_7_0_755_inst : InterlockBuffer generic map ( -- 
        name => "W_index2_755_delayed_7_0_755_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => index2_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => index2_755_delayed_7_0_757,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_437_inst
    process(sliced_v11_309) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v11_309(7 downto 0);
      a11_438 <= tmp_var; -- 
    end process;
    -- interlock type_cast_441_inst
    process(sliced_v12_313) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v12_313(7 downto 0);
      a12_442 <= tmp_var; -- 
    end process;
    -- interlock type_cast_445_inst
    process(sliced_v13_317) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v13_317(7 downto 0);
      a13_446 <= tmp_var; -- 
    end process;
    -- interlock type_cast_449_inst
    process(sliced_v14_321) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v14_321(7 downto 0);
      a14_450 <= tmp_var; -- 
    end process;
    -- interlock type_cast_453_inst
    process(sliced_v15_325) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v15_325(7 downto 0);
      a15_454 <= tmp_var; -- 
    end process;
    -- interlock type_cast_457_inst
    process(sliced_v16_329) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v16_329(7 downto 0);
      a16_458 <= tmp_var; -- 
    end process;
    -- interlock type_cast_461_inst
    process(sliced_v17_333) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v17_333(7 downto 0);
      a17_462 <= tmp_var; -- 
    end process;
    -- interlock type_cast_465_inst
    process(sliced_v18_337) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v18_337(7 downto 0);
      a18_466 <= tmp_var; -- 
    end process;
    -- interlock type_cast_469_inst
    process(sliced_v21_341) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v21_341(7 downto 0);
      a21_470 <= tmp_var; -- 
    end process;
    -- interlock type_cast_473_inst
    process(sliced_v22_345) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v22_345(7 downto 0);
      a22_474 <= tmp_var; -- 
    end process;
    -- interlock type_cast_477_inst
    process(sliced_v23_349) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v23_349(7 downto 0);
      a23_478 <= tmp_var; -- 
    end process;
    -- interlock type_cast_481_inst
    process(sliced_v24_353) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v24_353(7 downto 0);
      a24_482 <= tmp_var; -- 
    end process;
    -- interlock type_cast_485_inst
    process(sliced_v25_357) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v25_357(7 downto 0);
      a25_486 <= tmp_var; -- 
    end process;
    -- interlock type_cast_489_inst
    process(sliced_v26_361) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v26_361(7 downto 0);
      a26_490 <= tmp_var; -- 
    end process;
    -- interlock type_cast_493_inst
    process(sliced_v27_365) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v27_365(7 downto 0);
      a27_494 <= tmp_var; -- 
    end process;
    -- interlock type_cast_497_inst
    process(sliced_v28_369) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v28_369(7 downto 0);
      a28_498 <= tmp_var; -- 
    end process;
    -- interlock type_cast_501_inst
    process(sliced_v31_373) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v31_373(7 downto 0);
      a31_502 <= tmp_var; -- 
    end process;
    -- interlock type_cast_505_inst
    process(sliced_v32_377) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v32_377(7 downto 0);
      a32_506 <= tmp_var; -- 
    end process;
    -- interlock type_cast_509_inst
    process(sliced_v33_381) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v33_381(7 downto 0);
      a33_510 <= tmp_var; -- 
    end process;
    -- interlock type_cast_513_inst
    process(sliced_v34_385) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v34_385(7 downto 0);
      a34_514 <= tmp_var; -- 
    end process;
    -- interlock type_cast_517_inst
    process(sliced_v35_389) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v35_389(7 downto 0);
      a35_518 <= tmp_var; -- 
    end process;
    -- interlock type_cast_521_inst
    process(sliced_v36_393) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v36_393(7 downto 0);
      a36_522 <= tmp_var; -- 
    end process;
    -- interlock type_cast_525_inst
    process(sliced_v37_397) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v37_397(7 downto 0);
      a37_526 <= tmp_var; -- 
    end process;
    -- interlock type_cast_529_inst
    process(sliced_v38_401) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v38_401(7 downto 0);
      a38_530 <= tmp_var; -- 
    end process;
    -- interlock type_cast_533_inst
    process(sliced_v41_405) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v41_405(7 downto 0);
      a41_534 <= tmp_var; -- 
    end process;
    -- interlock type_cast_537_inst
    process(sliced_v42_409) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v42_409(7 downto 0);
      a42_538 <= tmp_var; -- 
    end process;
    -- interlock type_cast_541_inst
    process(sliced_v43_413) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v43_413(7 downto 0);
      a43_542 <= tmp_var; -- 
    end process;
    -- interlock type_cast_545_inst
    process(sliced_v44_417) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v44_417(7 downto 0);
      a44_546 <= tmp_var; -- 
    end process;
    -- interlock type_cast_549_inst
    process(sliced_v45_421) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v45_421(7 downto 0);
      a45_550 <= tmp_var; -- 
    end process;
    -- interlock type_cast_553_inst
    process(sliced_v46_425) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v46_425(7 downto 0);
      a46_554 <= tmp_var; -- 
    end process;
    -- interlock type_cast_557_inst
    process(sliced_v47_429) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v47_429(7 downto 0);
      a47_558 <= tmp_var; -- 
    end process;
    -- interlock type_cast_561_inst
    process(sliced_v48_433) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := sliced_v48_433(7 downto 0);
      a48_562 <= tmp_var; -- 
    end process;
    -- interlock type_cast_764_inst
    process(out1_586) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := out1_586(7 downto 0);
      type_cast_764_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_766_inst
    process(out2_610) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := out2_610(7 downto 0);
      type_cast_766_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_770_inst
    process(out3_634) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := out3_634(7 downto 0);
      type_cast_770_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_772_inst
    process(out4_658) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := out4_658(7 downto 0);
      type_cast_772_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_776_inst
    process(out5_682) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := out5_682(7 downto 0);
      type_cast_776_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_778_inst
    process(out6_706) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := out6_706(7 downto 0);
      type_cast_778_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_781_inst
    process(out7_730) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := out7_730(7 downto 0);
      type_cast_781_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_783_inst
    process(out8_754) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := out8_754(7 downto 0);
      type_cast_783_wire <= tmp_var; -- 
    end process;
    type_cast_791_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_791_inst_req_0;
      type_cast_791_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_791_inst_req_1;
      type_cast_791_inst_ack_1<= rack(0);
      type_cast_791_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_791_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => out1_586,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- binary operator CONCAT_u16_u32_774_inst
    process(CONCAT_u8_u16_767_wire, CONCAT_u8_u16_773_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_767_wire, CONCAT_u8_u16_773_wire, tmp_var);
      CONCAT_u16_u32_774_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_785_inst
    process(CONCAT_u8_u16_779_wire, CONCAT_u8_u16_784_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_779_wire, CONCAT_u8_u16_784_wire, tmp_var);
      CONCAT_u16_u32_785_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u64_786_inst
    process(CONCAT_u16_u32_774_wire, CONCAT_u16_u32_785_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u16_u32_774_wire, CONCAT_u16_u32_785_wire, tmp_var);
      CONCAT_u32_u64_786_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_767_inst
    process(type_cast_764_wire, type_cast_766_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_764_wire, type_cast_766_wire, tmp_var);
      CONCAT_u8_u16_767_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_773_inst
    process(type_cast_770_wire, type_cast_772_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_770_wire, type_cast_772_wire, tmp_var);
      CONCAT_u8_u16_773_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_779_inst
    process(type_cast_776_wire, type_cast_778_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_776_wire, type_cast_778_wire, tmp_var);
      CONCAT_u8_u16_779_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_784_inst
    process(type_cast_781_wire, type_cast_783_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_781_wire, type_cast_783_wire, tmp_var);
      CONCAT_u8_u16_784_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_566_inst
    process(a11_438, a21_470) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a11_438, a21_470, tmp_var);
      SGT_i8_u1_566_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_574_inst
    process(a31_502, a41_534) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a31_502, a41_534, tmp_var);
      SGT_i8_u1_574_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_582_inst
    process(t11_570, t12_578) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t11_570, t12_578, tmp_var);
      SGT_i8_u1_582_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_590_inst
    process(a12_442, a22_474) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a12_442, a22_474, tmp_var);
      SGT_i8_u1_590_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_598_inst
    process(a32_506, a42_538) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a32_506, a42_538, tmp_var);
      SGT_i8_u1_598_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_606_inst
    process(t21_594, t22_602) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t21_594, t22_602, tmp_var);
      SGT_i8_u1_606_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_614_inst
    process(a13_446, a23_478) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a13_446, a23_478, tmp_var);
      SGT_i8_u1_614_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_622_inst
    process(a33_510, a43_542) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a33_510, a43_542, tmp_var);
      SGT_i8_u1_622_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_630_inst
    process(t31_618, t32_626) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t31_618, t32_626, tmp_var);
      SGT_i8_u1_630_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_638_inst
    process(a14_450, a24_482) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a14_450, a24_482, tmp_var);
      SGT_i8_u1_638_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_646_inst
    process(a34_514, a44_546) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a34_514, a44_546, tmp_var);
      SGT_i8_u1_646_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_654_inst
    process(t41_642, t42_650) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t41_642, t42_650, tmp_var);
      SGT_i8_u1_654_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_662_inst
    process(a15_454, a25_486) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a15_454, a25_486, tmp_var);
      SGT_i8_u1_662_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_670_inst
    process(a35_518, a45_550) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a35_518, a45_550, tmp_var);
      SGT_i8_u1_670_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_678_inst
    process(t51_666, t52_674) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t51_666, t52_674, tmp_var);
      SGT_i8_u1_678_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_686_inst
    process(a16_458, a26_490) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a16_458, a26_490, tmp_var);
      SGT_i8_u1_686_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_694_inst
    process(a36_522, a46_554) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a36_522, a46_554, tmp_var);
      SGT_i8_u1_694_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_702_inst
    process(t61_690, t62_698) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t61_690, t62_698, tmp_var);
      SGT_i8_u1_702_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_710_inst
    process(a17_462, a27_494) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a17_462, a27_494, tmp_var);
      SGT_i8_u1_710_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_718_inst
    process(a37_526, a47_558) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a37_526, a47_558, tmp_var);
      SGT_i8_u1_718_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_726_inst
    process(t71_714, t72_722) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t71_714, t72_722, tmp_var);
      SGT_i8_u1_726_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_734_inst
    process(a18_466, a28_498) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a18_466, a28_498, tmp_var);
      SGT_i8_u1_734_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_742_inst
    process(a38_530, a48_562) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a38_530, a48_562, tmp_var);
      SGT_i8_u1_742_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i8_u1_750_inst
    process(t81_738, t82_746) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t81_738, t82_746, tmp_var);
      SGT_i8_u1_750_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_297_call call_stmt_293_call call_stmt_301_call call_stmt_305_call 
    readModule_maxPool_call_group_0: Block -- 
      signal data_in: std_logic_vector(159 downto 0);
      signal data_out: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 6, 1 => 6, 2 => 6, 3 => 6);
      -- 
    begin -- 
      reqL_unguarded(3) <= call_stmt_297_call_req_0;
      reqL_unguarded(2) <= call_stmt_293_call_req_0;
      reqL_unguarded(1) <= call_stmt_301_call_req_0;
      reqL_unguarded(0) <= call_stmt_305_call_req_0;
      call_stmt_297_call_ack_0 <= ackL_unguarded(3);
      call_stmt_293_call_ack_0 <= ackL_unguarded(2);
      call_stmt_301_call_ack_0 <= ackL_unguarded(1);
      call_stmt_305_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= call_stmt_297_call_req_1;
      reqR_unguarded(2) <= call_stmt_293_call_req_1;
      reqR_unguarded(1) <= call_stmt_301_call_req_1;
      reqR_unguarded(0) <= call_stmt_305_call_req_1;
      call_stmt_297_call_ack_1 <= ackR_unguarded(3);
      call_stmt_293_call_ack_1 <= ackR_unguarded(2);
      call_stmt_301_call_ack_1 <= ackR_unguarded(1);
      call_stmt_305_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      readModule_maxPool_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "readModule_maxPool_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      readModule_maxPool_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "readModule_maxPool_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      readModule_maxPool_call_group_0_accessRegulator_2: access_regulator_base generic map (name => "readModule_maxPool_call_group_0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      readModule_maxPool_call_group_0_accessRegulator_3: access_regulator_base generic map (name => "readModule_maxPool_call_group_0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      readModule_maxPool_call_group_0_gI: SplitGuardInterface generic map(name => "readModule_maxPool_call_group_0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= index1_buffer & addr2_buffer & index1_buffer & addr1_buffer & index1_buffer & addr3_buffer & index1_buffer & addr4_buffer;
      c2_297 <= data_out(255 downto 192);
      c1_293 <= data_out(191 downto 128);
      c3_301 <= data_out(127 downto 64);
      c4_305 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 160,
        owidth => 40,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 3,
        nreqs => 4,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => readModule_maxPool_call_reqs(0),
          ackR => readModule_maxPool_call_acks(0),
          dataR => readModule_maxPool_call_data(39 downto 0),
          tagR => readModule_maxPool_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 256,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 4) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => readModule_maxPool_return_acks(0), -- cross-over
          ackL => readModule_maxPool_return_reqs(0), -- cross-over
          dataL => readModule_maxPool_return_data(63 downto 0),
          tagL => readModule_maxPool_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_788_call 
    writeModule_maxPool_call_group_1: Block -- 
      signal data_in: std_logic_vector(103 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_788_call_req_0;
      call_stmt_788_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_788_call_req_1;
      call_stmt_788_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writeModule_maxPool_call_group_1_gI: SplitGuardInterface generic map(name => "writeModule_maxPool_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= index2_755_delayed_7_0_757 & addr_756_delayed_7_0_760 & CONCAT_u32_u64_786_wire;
      d1_788 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 104,
        owidth => 104,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writeModule_maxPool_call_reqs(0),
          ackR => writeModule_maxPool_call_acks(0),
          dataR => writeModule_maxPool_call_data(103 downto 0),
          tagR => writeModule_maxPool_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => writeModule_maxPool_return_acks(0), -- cross-over
          ackL => writeModule_maxPool_return_reqs(0), -- cross-over
          dataL => writeModule_maxPool_return_data(0 downto 0),
          tagL => writeModule_maxPool_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end maxPool4_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity memoryModule is -- 
  generic (tag_length : integer); 
  port ( -- 
    r_wbar : in  std_logic_vector(0 downto 0);
    addr : in  std_logic_vector(31 downto 0);
    data_in : in  std_logic_vector(63 downto 0);
    data_out : out  std_logic_vector(63 downto 0);
    MAIN_MEM_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
    MAIN_MEM_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    MAIN_MEM_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
    MAIN_MEM_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
    MAIN_MEM_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
    MAIN_MEM_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity memoryModule;
architecture memoryModule_arch of memoryModule is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 97)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal r_wbar_buffer :  std_logic_vector(0 downto 0);
  signal r_wbar_update_enable: Boolean;
  signal addr_buffer :  std_logic_vector(31 downto 0);
  signal addr_update_enable: Boolean;
  signal data_in_buffer :  std_logic_vector(63 downto 0);
  signal data_in_update_enable: Boolean;
  -- output port buffer signals
  signal data_out_buffer :  std_logic_vector(63 downto 0);
  signal data_out_update_enable: Boolean;
  signal memoryModule_CP_0_start: Boolean;
  signal memoryModule_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal CONCAT_u10_u110_50_inst_req_0 : boolean;
  signal CONCAT_u10_u110_50_inst_ack_0 : boolean;
  signal CONCAT_u10_u110_50_inst_req_1 : boolean;
  signal CONCAT_u10_u110_50_inst_ack_1 : boolean;
  signal WPIPE_MAIN_MEM_REQUEST_35_inst_req_0 : boolean;
  signal WPIPE_MAIN_MEM_REQUEST_35_inst_ack_0 : boolean;
  signal WPIPE_MAIN_MEM_REQUEST_35_inst_req_1 : boolean;
  signal WPIPE_MAIN_MEM_REQUEST_35_inst_ack_1 : boolean;
  signal RPIPE_MAIN_MEM_RESPONSE_53_inst_req_0 : boolean;
  signal RPIPE_MAIN_MEM_RESPONSE_53_inst_ack_0 : boolean;
  signal RPIPE_MAIN_MEM_RESPONSE_53_inst_req_1 : boolean;
  signal RPIPE_MAIN_MEM_RESPONSE_53_inst_ack_1 : boolean;
  signal slice_54_inst_req_0 : boolean;
  signal slice_54_inst_ack_0 : boolean;
  signal slice_54_inst_req_1 : boolean;
  signal slice_54_inst_ack_1 : boolean;
  signal RPIPE_MAIN_MEM_RESPONSE_57_inst_req_0 : boolean;
  signal RPIPE_MAIN_MEM_RESPONSE_57_inst_ack_0 : boolean;
  signal RPIPE_MAIN_MEM_RESPONSE_57_inst_req_1 : boolean;
  signal RPIPE_MAIN_MEM_RESPONSE_57_inst_ack_1 : boolean;
  signal slice_58_inst_req_0 : boolean;
  signal slice_58_inst_ack_0 : boolean;
  signal slice_58_inst_req_1 : boolean;
  signal slice_58_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "memoryModule_input_buffer", -- 
      buffer_size => 2,
      bypass_flag => false,
      data_width => tag_length + 97) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= r_wbar;
  r_wbar_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(32 downto 1) <= addr;
  addr_buffer <= in_buffer_data_out(32 downto 1);
  in_buffer_data_in(96 downto 33) <= data_in;
  data_in_buffer <= in_buffer_data_out(96 downto 33);
  in_buffer_data_in(tag_length + 96 downto 97) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 96 downto 97);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 15);
    constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 15);
    constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 5); -- 
  begin -- 
    preds <= r_wbar_update_enable & addr_update_enable & data_in_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  memoryModule_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "memoryModule_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= data_out_buffer;
  data_out <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 15);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= memoryModule_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  data_out_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 27) := "data_out_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_data_out_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => data_out_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 15,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= memoryModule_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= memoryModule_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  memoryModule_CP_0: Block -- control-path 
    signal memoryModule_CP_0_elements: BooleanArray(34 downto 0);
    -- 
  begin -- 
    memoryModule_CP_0_elements(0) <= memoryModule_CP_0_start;
    memoryModule_CP_0_symbol <= memoryModule_CP_0_elements(34);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	6 
    -- CP-element group 1: 	15 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 assign_stmt_51_to_assign_stmt_59/$entry
      -- 
    memoryModule_CP_0_elements(1) <= memoryModule_CP_0_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	8 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	30 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_51_to_assign_stmt_59/r_wbar_update_enable
      -- CP-element group 2: 	 assign_stmt_51_to_assign_stmt_59/r_wbar_update_enable_out
      -- 
    memoryModule_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "memoryModule_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= memoryModule_CP_0_elements(8);
      gj_memoryModule_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryModule_CP_0_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	8 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	31 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_51_to_assign_stmt_59/addr_update_enable
      -- CP-element group 3: 	 assign_stmt_51_to_assign_stmt_59/addr_update_enable_out
      -- 
    memoryModule_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "memoryModule_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= memoryModule_CP_0_elements(8);
      gj_memoryModule_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryModule_CP_0_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	8 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	32 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_51_to_assign_stmt_59/data_in_update_enable_out
      -- CP-element group 4: 	 assign_stmt_51_to_assign_stmt_59/data_in_update_enable
      -- 
    memoryModule_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "memoryModule_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= memoryModule_CP_0_elements(8);
      gj_memoryModule_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryModule_CP_0_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	33 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	22 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_51_to_assign_stmt_59/data_out_update_enable
      -- CP-element group 5: 	 assign_stmt_51_to_assign_stmt_59/data_out_update_enable_in
      -- 
    memoryModule_CP_0_elements(5) <= memoryModule_CP_0_elements(33);
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	1 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	8 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_51_to_assign_stmt_59/CONCAT_u10_u110_50_sample_start_
      -- CP-element group 6: 	 assign_stmt_51_to_assign_stmt_59/CONCAT_u10_u110_50_Sample/$entry
      -- CP-element group 6: 	 assign_stmt_51_to_assign_stmt_59/CONCAT_u10_u110_50_Sample/rr
      -- 
    rr_21_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_21_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memoryModule_CP_0_elements(6), ack => CONCAT_u10_u110_50_inst_req_0); -- 
    memoryModule_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "memoryModule_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memoryModule_CP_0_elements(1) & memoryModule_CP_0_elements(8);
      gj_memoryModule_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryModule_CP_0_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: marked-predecessors 
    -- CP-element group 7: 	9 
    -- CP-element group 7: 	11 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	9 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_51_to_assign_stmt_59/CONCAT_u10_u110_50_update_start_
      -- CP-element group 7: 	 assign_stmt_51_to_assign_stmt_59/CONCAT_u10_u110_50_Update/$entry
      -- CP-element group 7: 	 assign_stmt_51_to_assign_stmt_59/CONCAT_u10_u110_50_Update/cr
      -- 
    cr_26_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_26_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memoryModule_CP_0_elements(7), ack => CONCAT_u10_u110_50_inst_req_1); -- 
    memoryModule_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "memoryModule_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memoryModule_CP_0_elements(9) & memoryModule_CP_0_elements(11);
      gj_memoryModule_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryModule_CP_0_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: 	3 
    -- CP-element group 8: 	4 
    -- CP-element group 8: 	6 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_51_to_assign_stmt_59/CONCAT_u10_u110_50_sample_completed_
      -- CP-element group 8: 	 assign_stmt_51_to_assign_stmt_59/CONCAT_u10_u110_50_Sample/$exit
      -- CP-element group 8: 	 assign_stmt_51_to_assign_stmt_59/CONCAT_u10_u110_50_Sample/ra
      -- 
    ra_22_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u10_u110_50_inst_ack_0, ack => memoryModule_CP_0_elements(8)); -- 
    -- CP-element group 9:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	7 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: marked-successors 
    -- CP-element group 9: 	7 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_51_to_assign_stmt_59/CONCAT_u10_u110_50_update_completed_
      -- CP-element group 9: 	 assign_stmt_51_to_assign_stmt_59/CONCAT_u10_u110_50_Update/$exit
      -- CP-element group 9: 	 assign_stmt_51_to_assign_stmt_59/CONCAT_u10_u110_50_Update/ca
      -- 
    ca_27_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u10_u110_50_inst_ack_1, ack => memoryModule_CP_0_elements(9)); -- 
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_51_to_assign_stmt_59/WPIPE_MAIN_MEM_REQUEST_35_sample_start_
      -- CP-element group 10: 	 assign_stmt_51_to_assign_stmt_59/WPIPE_MAIN_MEM_REQUEST_35_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_51_to_assign_stmt_59/WPIPE_MAIN_MEM_REQUEST_35_Sample/req
      -- 
    req_35_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_35_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memoryModule_CP_0_elements(10), ack => WPIPE_MAIN_MEM_REQUEST_35_inst_req_0); -- 
    memoryModule_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "memoryModule_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memoryModule_CP_0_elements(9) & memoryModule_CP_0_elements(12);
      gj_memoryModule_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryModule_CP_0_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	7 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 assign_stmt_51_to_assign_stmt_59/WPIPE_MAIN_MEM_REQUEST_35_sample_completed_
      -- CP-element group 11: 	 assign_stmt_51_to_assign_stmt_59/WPIPE_MAIN_MEM_REQUEST_35_update_start_
      -- CP-element group 11: 	 assign_stmt_51_to_assign_stmt_59/WPIPE_MAIN_MEM_REQUEST_35_Sample/$exit
      -- CP-element group 11: 	 assign_stmt_51_to_assign_stmt_59/WPIPE_MAIN_MEM_REQUEST_35_Sample/ack
      -- CP-element group 11: 	 assign_stmt_51_to_assign_stmt_59/WPIPE_MAIN_MEM_REQUEST_35_Update/$entry
      -- CP-element group 11: 	 assign_stmt_51_to_assign_stmt_59/WPIPE_MAIN_MEM_REQUEST_35_Update/req
      -- 
    ack_36_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_MAIN_MEM_REQUEST_35_inst_ack_0, ack => memoryModule_CP_0_elements(11)); -- 
    req_40_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_40_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memoryModule_CP_0_elements(11), ack => WPIPE_MAIN_MEM_REQUEST_35_inst_req_1); -- 
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	29 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_51_to_assign_stmt_59/WPIPE_MAIN_MEM_REQUEST_35_update_completed_
      -- CP-element group 12: 	 assign_stmt_51_to_assign_stmt_59/WPIPE_MAIN_MEM_REQUEST_35_Update/$exit
      -- CP-element group 12: 	 assign_stmt_51_to_assign_stmt_59/WPIPE_MAIN_MEM_REQUEST_35_Update/ack
      -- 
    ack_41_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_MAIN_MEM_REQUEST_35_inst_ack_1, ack => memoryModule_CP_0_elements(12)); -- 
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	18 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	19 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	19 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_51_to_assign_stmt_59/slice_54_sample_start_
      -- CP-element group 13: 	 assign_stmt_51_to_assign_stmt_59/slice_54_Sample/$entry
      -- CP-element group 13: 	 assign_stmt_51_to_assign_stmt_59/slice_54_Sample/rr
      -- 
    rr_63_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_63_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memoryModule_CP_0_elements(13), ack => slice_54_inst_req_0); -- 
    memoryModule_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "memoryModule_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memoryModule_CP_0_elements(18) & memoryModule_CP_0_elements(19);
      gj_memoryModule_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryModule_CP_0_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	20 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	20 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_51_to_assign_stmt_59/slice_54_update_start_
      -- CP-element group 14: 	 assign_stmt_51_to_assign_stmt_59/slice_54_Update/$entry
      -- CP-element group 14: 	 assign_stmt_51_to_assign_stmt_59/slice_54_Update/cr
      -- 
    cr_68_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_68_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memoryModule_CP_0_elements(14), ack => slice_54_inst_req_1); -- 
    memoryModule_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "memoryModule_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= memoryModule_CP_0_elements(20);
      gj_memoryModule_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryModule_CP_0_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	1 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	18 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_53_sample_start_
      -- CP-element group 15: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_53_Sample/$entry
      -- CP-element group 15: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_53_Sample/rr
      -- 
    rr_53_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_53_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memoryModule_CP_0_elements(15), ack => RPIPE_MAIN_MEM_RESPONSE_53_inst_req_0); -- 
    memoryModule_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "memoryModule_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memoryModule_CP_0_elements(1) & memoryModule_CP_0_elements(18);
      gj_memoryModule_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryModule_CP_0_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	17 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	19 
    -- CP-element group 16: 	26 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_53_update_start_
      -- CP-element group 16: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_53_Update/$entry
      -- CP-element group 16: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_53_Update/cr
      -- 
    cr_58_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_58_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memoryModule_CP_0_elements(16), ack => RPIPE_MAIN_MEM_RESPONSE_53_inst_req_1); -- 
    memoryModule_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "memoryModule_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= memoryModule_CP_0_elements(17) & memoryModule_CP_0_elements(19) & memoryModule_CP_0_elements(26);
      gj_memoryModule_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryModule_CP_0_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	16 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_53_sample_completed_
      -- CP-element group 17: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_53_Sample/$exit
      -- CP-element group 17: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_53_Sample/ra
      -- 
    ra_54_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_MAIN_MEM_RESPONSE_53_inst_ack_0, ack => memoryModule_CP_0_elements(17)); -- 
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	13 
    -- CP-element group 18: 	23 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	15 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_53_update_completed_
      -- CP-element group 18: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_53_Update/$exit
      -- CP-element group 18: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_53_Update/ca
      -- 
    ca_59_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_MAIN_MEM_RESPONSE_53_inst_ack_1, ack => memoryModule_CP_0_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: 	16 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 assign_stmt_51_to_assign_stmt_59/slice_54_sample_completed_
      -- CP-element group 19: 	 assign_stmt_51_to_assign_stmt_59/slice_54_Sample/$exit
      -- CP-element group 19: 	 assign_stmt_51_to_assign_stmt_59/slice_54_Sample/ra
      -- 
    ra_64_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_54_inst_ack_0, ack => memoryModule_CP_0_elements(19)); -- 
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	29 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	14 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 assign_stmt_51_to_assign_stmt_59/slice_54_update_completed_
      -- CP-element group 20: 	 assign_stmt_51_to_assign_stmt_59/slice_54_Update/$exit
      -- CP-element group 20: 	 assign_stmt_51_to_assign_stmt_59/slice_54_Update/ca
      -- 
    ca_69_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_54_inst_ack_1, ack => memoryModule_CP_0_elements(20)); -- 
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	26 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	27 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	27 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 assign_stmt_51_to_assign_stmt_59/slice_58_sample_start_
      -- CP-element group 21: 	 assign_stmt_51_to_assign_stmt_59/slice_58_Sample/$entry
      -- CP-element group 21: 	 assign_stmt_51_to_assign_stmt_59/slice_58_Sample/rr
      -- 
    rr_91_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_91_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memoryModule_CP_0_elements(21), ack => slice_58_inst_req_0); -- 
    memoryModule_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "memoryModule_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memoryModule_CP_0_elements(26) & memoryModule_CP_0_elements(27);
      gj_memoryModule_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryModule_CP_0_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	5 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	28 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	28 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 assign_stmt_51_to_assign_stmt_59/slice_58_update_start_
      -- CP-element group 22: 	 assign_stmt_51_to_assign_stmt_59/slice_58_Update/$entry
      -- CP-element group 22: 	 assign_stmt_51_to_assign_stmt_59/slice_58_Update/cr
      -- 
    cr_96_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_96_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memoryModule_CP_0_elements(22), ack => slice_58_inst_req_1); -- 
    memoryModule_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "memoryModule_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memoryModule_CP_0_elements(5) & memoryModule_CP_0_elements(28);
      gj_memoryModule_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryModule_CP_0_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	18 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	26 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_57_sample_start_
      -- CP-element group 23: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_57_Sample/$entry
      -- CP-element group 23: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_57_Sample/rr
      -- 
    rr_81_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_81_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memoryModule_CP_0_elements(23), ack => RPIPE_MAIN_MEM_RESPONSE_57_inst_req_0); -- 
    memoryModule_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "memoryModule_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memoryModule_CP_0_elements(18) & memoryModule_CP_0_elements(26);
      gj_memoryModule_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryModule_CP_0_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	25 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	27 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_57_update_start_
      -- CP-element group 24: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_57_Update/$entry
      -- CP-element group 24: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_57_Update/cr
      -- 
    cr_86_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_86_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memoryModule_CP_0_elements(24), ack => RPIPE_MAIN_MEM_RESPONSE_57_inst_req_1); -- 
    memoryModule_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "memoryModule_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memoryModule_CP_0_elements(25) & memoryModule_CP_0_elements(27);
      gj_memoryModule_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryModule_CP_0_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	24 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_57_sample_completed_
      -- CP-element group 25: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_57_Sample/$exit
      -- CP-element group 25: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_57_Sample/ra
      -- 
    ra_82_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_MAIN_MEM_RESPONSE_57_inst_ack_0, ack => memoryModule_CP_0_elements(25)); -- 
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	21 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	16 
    -- CP-element group 26: 	23 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_57_update_completed_
      -- CP-element group 26: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_57_Update/$exit
      -- CP-element group 26: 	 assign_stmt_51_to_assign_stmt_59/RPIPE_MAIN_MEM_RESPONSE_57_Update/ca
      -- 
    ca_87_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_MAIN_MEM_RESPONSE_57_inst_ack_1, ack => memoryModule_CP_0_elements(26)); -- 
    -- CP-element group 27:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	21 
    -- CP-element group 27: successors 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	21 
    -- CP-element group 27: 	24 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_51_to_assign_stmt_59/slice_58_sample_completed_
      -- CP-element group 27: 	 assign_stmt_51_to_assign_stmt_59/slice_58_Sample/$exit
      -- CP-element group 27: 	 assign_stmt_51_to_assign_stmt_59/slice_58_Sample/ra
      -- 
    ra_92_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_58_inst_ack_0, ack => memoryModule_CP_0_elements(27)); -- 
    -- CP-element group 28:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	22 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	22 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 assign_stmt_51_to_assign_stmt_59/slice_58_update_completed_
      -- CP-element group 28: 	 assign_stmt_51_to_assign_stmt_59/slice_58_Update/$exit
      -- CP-element group 28: 	 assign_stmt_51_to_assign_stmt_59/slice_58_Update/ca
      -- 
    ca_97_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_58_inst_ack_1, ack => memoryModule_CP_0_elements(28)); -- 
    -- CP-element group 29:  join  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	12 
    -- CP-element group 29: 	20 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	34 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 assign_stmt_51_to_assign_stmt_59/$exit
      -- 
    memoryModule_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "memoryModule_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= memoryModule_CP_0_elements(12) & memoryModule_CP_0_elements(20) & memoryModule_CP_0_elements(28);
      gj_memoryModule_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryModule_CP_0_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  place  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	2 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 r_wbar_update_enable
      -- 
    memoryModule_CP_0_elements(30) <= memoryModule_CP_0_elements(2);
    -- CP-element group 31:  place  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	3 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 addr_update_enable
      -- 
    memoryModule_CP_0_elements(31) <= memoryModule_CP_0_elements(3);
    -- CP-element group 32:  place  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	4 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 data_in_update_enable
      -- 
    memoryModule_CP_0_elements(32) <= memoryModule_CP_0_elements(4);
    -- CP-element group 33:  place  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	5 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 data_out_update_enable
      -- 
    -- CP-element group 34:  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	29 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 $exit
      -- 
    memoryModule_CP_0_elements(34) <= memoryModule_CP_0_elements(29);
    --  hookup: inputs to control-path 
    memoryModule_CP_0_elements(33) <= data_out_update_enable;
    -- hookup: output from control-path 
    r_wbar_update_enable <= memoryModule_CP_0_elements(30);
    addr_update_enable <= memoryModule_CP_0_elements(31);
    data_in_update_enable <= memoryModule_CP_0_elements(32);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u10_u110_50_wire : std_logic_vector(109 downto 0);
    signal CONCAT_u1_u2_39_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u2_u10_42_wire : std_logic_vector(9 downto 0);
    signal CONCAT_u36_u100_49_wire : std_logic_vector(99 downto 0);
    signal CONCAT_u4_u36_47_wire : std_logic_vector(35 downto 0);
    signal RPIPE_MAIN_MEM_RESPONSE_53_wire : std_logic_vector(64 downto 0);
    signal RPIPE_MAIN_MEM_RESPONSE_57_wire : std_logic_vector(64 downto 0);
    signal error_55 : std_logic_vector(0 downto 0);
    signal type_cast_37_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_41_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_45_wire_constant : std_logic_vector(3 downto 0);
    -- 
  begin -- 
    type_cast_37_wire_constant <= "0";
    type_cast_41_wire_constant <= "00000001";
    type_cast_45_wire_constant <= "0000";
    slice_54_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_54_inst_req_0;
      slice_54_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_54_inst_req_1;
      slice_54_inst_ack_1<= update_ack(0);
      slice_54_inst: SliceSplitProtocol generic map(name => "slice_54_inst", in_data_width => 65, high_index => 64, low_index => 64, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => RPIPE_MAIN_MEM_RESPONSE_53_wire, dout => error_55, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_58_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_58_inst_req_0;
      slice_58_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_58_inst_req_1;
      slice_58_inst_ack_1<= update_ack(0);
      slice_58_inst: SliceSplitProtocol generic map(name => "slice_58_inst", in_data_width => 65, high_index => 63, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => RPIPE_MAIN_MEM_RESPONSE_57_wire, dout => data_out_buffer, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- shared split operator group (0) : CONCAT_u10_u110_50_inst 
    ApConcat_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(109 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u2_u10_42_wire & CONCAT_u36_u100_49_wire;
      CONCAT_u10_u110_50_wire <= data_out(109 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u10_u110_50_inst_req_0;
      CONCAT_u10_u110_50_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u10_u110_50_inst_req_1;
      CONCAT_u10_u110_50_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_0_gI: SplitGuardInterface generic map(name => "ApConcat_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 10,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 100, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 110,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator CONCAT_u1_u2_39_inst
    process(type_cast_37_wire_constant, r_wbar_buffer) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_37_wire_constant, r_wbar_buffer, tmp_var);
      CONCAT_u1_u2_39_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u10_42_inst
    process(CONCAT_u1_u2_39_wire) -- 
      variable tmp_var : std_logic_vector(9 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_39_wire, type_cast_41_wire_constant, tmp_var);
      CONCAT_u2_u10_42_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u36_u100_49_inst
    process(CONCAT_u4_u36_47_wire, data_in_buffer) -- 
      variable tmp_var : std_logic_vector(99 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u4_u36_47_wire, data_in_buffer, tmp_var);
      CONCAT_u36_u100_49_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u36_47_inst
    process(type_cast_45_wire_constant, addr_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_45_wire_constant, addr_buffer, tmp_var);
      CONCAT_u4_u36_47_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_MAIN_MEM_RESPONSE_57_inst RPIPE_MAIN_MEM_RESPONSE_53_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(129 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_MAIN_MEM_RESPONSE_57_inst_req_0;
      reqL_unguarded(0) <= RPIPE_MAIN_MEM_RESPONSE_53_inst_req_0;
      RPIPE_MAIN_MEM_RESPONSE_57_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_MAIN_MEM_RESPONSE_53_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_MAIN_MEM_RESPONSE_57_inst_req_1;
      reqR_unguarded(0) <= RPIPE_MAIN_MEM_RESPONSE_53_inst_req_1;
      RPIPE_MAIN_MEM_RESPONSE_57_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_MAIN_MEM_RESPONSE_53_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      RPIPE_MAIN_MEM_RESPONSE_57_wire <= data_out(129 downto 65);
      RPIPE_MAIN_MEM_RESPONSE_53_wire <= data_out(64 downto 0);
      MAIN_MEM_RESPONSE_read_0_gI: SplitGuardInterface generic map(name => "MAIN_MEM_RESPONSE_read_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      MAIN_MEM_RESPONSE_read_0: InputPortRevised -- 
        generic map ( name => "MAIN_MEM_RESPONSE_read_0", data_width => 65,  num_reqs => 2,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => MAIN_MEM_RESPONSE_pipe_read_req(0),
          oack => MAIN_MEM_RESPONSE_pipe_read_ack(0),
          odata => MAIN_MEM_RESPONSE_pipe_read_data(64 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_MAIN_MEM_REQUEST_35_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_MAIN_MEM_REQUEST_35_inst_req_0;
      WPIPE_MAIN_MEM_REQUEST_35_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_MAIN_MEM_REQUEST_35_inst_req_1;
      WPIPE_MAIN_MEM_REQUEST_35_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= CONCAT_u10_u110_50_wire;
      MAIN_MEM_REQUEST_write_0_gI: SplitGuardInterface generic map(name => "MAIN_MEM_REQUEST_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      MAIN_MEM_REQUEST_write_0: OutputPortRevised -- 
        generic map ( name => "MAIN_MEM_REQUEST", data_width => 110, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => MAIN_MEM_REQUEST_pipe_write_req(0),
          oack => MAIN_MEM_REQUEST_pipe_write_ack(0),
          odata => MAIN_MEM_REQUEST_pipe_write_data(109 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end memoryModule_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity readModule1 is -- 
  generic (tag_length : integer); 
  port ( -- 
    address : in  std_logic_vector(31 downto 0);
    data : out  std_logic_vector(63 downto 0);
    memoryModule_call_reqs : out  std_logic_vector(0 downto 0);
    memoryModule_call_acks : in   std_logic_vector(0 downto 0);
    memoryModule_call_data : out  std_logic_vector(96 downto 0);
    memoryModule_call_tag  :  out  std_logic_vector(0 downto 0);
    memoryModule_return_reqs : out  std_logic_vector(0 downto 0);
    memoryModule_return_acks : in   std_logic_vector(0 downto 0);
    memoryModule_return_data : in   std_logic_vector(63 downto 0);
    memoryModule_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity readModule1;
architecture readModule1_arch of readModule1 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal address_buffer :  std_logic_vector(31 downto 0);
  signal address_update_enable: Boolean;
  -- output port buffer signals
  signal data_buffer :  std_logic_vector(63 downto 0);
  signal data_update_enable: Boolean;
  signal readModule1_CP_1651_start: Boolean;
  signal readModule1_CP_1651_symbol: Boolean;
  -- volatile/operator module components. 
  component memoryModule is -- 
    generic (tag_length : integer); 
    port ( -- 
      r_wbar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(31 downto 0);
      data_in : in  std_logic_vector(63 downto 0);
      data_out : out  std_logic_vector(63 downto 0);
      MAIN_MEM_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MAIN_MEM_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MAIN_MEM_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      MAIN_MEM_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      MAIN_MEM_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      MAIN_MEM_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1042_call_req_0 : boolean;
  signal call_stmt_1042_call_ack_1 : boolean;
  signal call_stmt_1042_call_req_1 : boolean;
  signal call_stmt_1042_call_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "readModule1_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 32) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= address;
  address_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(tag_length + 31 downto 32) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 31 downto 32);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  readModule1_CP_1651_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "readModule1_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= data_buffer;
  data <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= readModule1_CP_1651_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= readModule1_CP_1651_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= readModule1_CP_1651_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  readModule1_CP_1651: Block -- control-path 
    signal readModule1_CP_1651_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    readModule1_CP_1651_elements(0) <= readModule1_CP_1651_start;
    readModule1_CP_1651_symbol <= readModule1_CP_1651_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_1042/call_stmt_1042_Sample/crr
      -- CP-element group 0: 	 call_stmt_1042/call_stmt_1042_update_start_
      -- CP-element group 0: 	 call_stmt_1042/call_stmt_1042_Sample/$entry
      -- CP-element group 0: 	 call_stmt_1042/$entry
      -- CP-element group 0: 	 call_stmt_1042/call_stmt_1042_sample_start_
      -- CP-element group 0: 	 call_stmt_1042/call_stmt_1042_Update/ccr
      -- CP-element group 0: 	 call_stmt_1042/call_stmt_1042_Update/$entry
      -- CP-element group 0: 	 $entry
      -- 
    crr_1664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_1651_elements(0), ack => call_stmt_1042_call_req_0); -- 
    ccr_1669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_1651_elements(0), ack => call_stmt_1042_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_1042/call_stmt_1042_sample_completed_
      -- CP-element group 1: 	 call_stmt_1042/call_stmt_1042_Sample/$exit
      -- CP-element group 1: 	 call_stmt_1042/call_stmt_1042_Sample/cra
      -- 
    cra_1665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1042_call_ack_0, ack => readModule1_CP_1651_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 call_stmt_1042/call_stmt_1042_update_completed_
      -- CP-element group 2: 	 call_stmt_1042/$exit
      -- CP-element group 2: 	 call_stmt_1042/call_stmt_1042_Update/cca
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_1042/call_stmt_1042_Update/$exit
      -- 
    cca_1670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1042_call_ack_1, ack => readModule1_CP_1651_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_1039_wire : std_logic_vector(31 downto 0);
    signal konst_1036_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1037_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1040_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_1036_wire_constant <= "1";
    konst_1037_wire_constant <= "00000000000000000000000000000000";
    konst_1040_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- binary operator ADD_u32_u32_1039_inst
    process(address_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address_buffer, konst_1037_wire_constant, tmp_var);
      ADD_u32_u32_1039_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_1042_call 
    memoryModule_call_group_0: Block -- 
      signal data_in: std_logic_vector(96 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1042_call_req_0;
      call_stmt_1042_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1042_call_req_1;
      call_stmt_1042_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      memoryModule_call_group_0_gI: SplitGuardInterface generic map(name => "memoryModule_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_1036_wire_constant & ADD_u32_u32_1039_wire & konst_1040_wire_constant;
      data_buffer <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 97,
        owidth => 97,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => memoryModule_call_reqs(0),
          ackR => memoryModule_call_acks(0),
          dataR => memoryModule_call_data(96 downto 0),
          tagR => memoryModule_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => memoryModule_return_acks(0), -- cross-over
          ackL => memoryModule_return_reqs(0), -- cross-over
          dataL => memoryModule_return_data(63 downto 0),
          tagL => memoryModule_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end readModule1_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity readModule_maxPool is -- 
  generic (tag_length : integer); 
  port ( -- 
    index : in  std_logic_vector(7 downto 0);
    address : in  std_logic_vector(31 downto 0);
    data : out  std_logic_vector(63 downto 0);
    memoryModule_call_reqs : out  std_logic_vector(0 downto 0);
    memoryModule_call_acks : in   std_logic_vector(0 downto 0);
    memoryModule_call_data : out  std_logic_vector(96 downto 0);
    memoryModule_call_tag  :  out  std_logic_vector(0 downto 0);
    memoryModule_return_reqs : out  std_logic_vector(0 downto 0);
    memoryModule_return_acks : in   std_logic_vector(0 downto 0);
    memoryModule_return_data : in   std_logic_vector(63 downto 0);
    memoryModule_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity readModule_maxPool;
architecture readModule_maxPool_arch of readModule_maxPool is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 40)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal index_buffer :  std_logic_vector(7 downto 0);
  signal index_update_enable: Boolean;
  signal address_buffer :  std_logic_vector(31 downto 0);
  signal address_update_enable: Boolean;
  -- output port buffer signals
  signal data_buffer :  std_logic_vector(63 downto 0);
  signal data_update_enable: Boolean;
  signal readModule_maxPool_CP_488_start: Boolean;
  signal readModule_maxPool_CP_488_symbol: Boolean;
  -- volatile/operator module components. 
  component memoryModule is -- 
    generic (tag_length : integer); 
    port ( -- 
      r_wbar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(31 downto 0);
      data_in : in  std_logic_vector(63 downto 0);
      data_out : out  std_logic_vector(63 downto 0);
      MAIN_MEM_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MAIN_MEM_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MAIN_MEM_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      MAIN_MEM_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      MAIN_MEM_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      MAIN_MEM_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_261_call_ack_1 : boolean;
  signal call_stmt_261_call_req_1 : boolean;
  signal call_stmt_261_call_ack_0 : boolean;
  signal call_stmt_261_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "readModule_maxPool_input_buffer", -- 
      buffer_size => 2,
      bypass_flag => false,
      data_width => tag_length + 40) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= index;
  index_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(39 downto 8) <= address;
  address_buffer <= in_buffer_data_out(39 downto 8);
  in_buffer_data_in(tag_length + 39 downto 40) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 39 downto 40);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 8);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 8);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= address_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  readModule_maxPool_CP_488_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "readModule_maxPool_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= data_buffer;
  data <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 8);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= readModule_maxPool_CP_488_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  data_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 23) := "data_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_data_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => data_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 8,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= readModule_maxPool_CP_488_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= readModule_maxPool_CP_488_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  readModule_maxPool_CP_488: Block -- control-path 
    signal readModule_maxPool_CP_488_elements: BooleanArray(12 downto 0);
    -- 
  begin -- 
    readModule_maxPool_CP_488_elements(0) <= readModule_maxPool_CP_488_start;
    readModule_maxPool_CP_488_symbol <= readModule_maxPool_CP_488_elements(12);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	5 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 call_stmt_261/$entry
      -- 
    readModule_maxPool_CP_488_elements(1) <= readModule_maxPool_CP_488_elements(0);
    -- CP-element group 2:  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	9 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 call_stmt_261/index_update_enable_out
      -- CP-element group 2: 	 call_stmt_261/index_update_enable
      -- 
    readModule_maxPool_CP_488_elements(2) <= false; 
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	7 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	10 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 call_stmt_261/address_update_enable_out
      -- CP-element group 3: 	 call_stmt_261/address_update_enable
      -- 
    readModule_maxPool_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 37) := "readModule_maxPool_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readModule_maxPool_CP_488_elements(7);
      gj_readModule_maxPool_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule_maxPool_CP_488_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	11 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	6 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 call_stmt_261/data_update_enable_in
      -- CP-element group 4: 	 call_stmt_261/data_update_enable
      -- 
    readModule_maxPool_CP_488_elements(4) <= readModule_maxPool_CP_488_elements(11);
    -- CP-element group 5:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	1 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	7 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_261/call_stmt_261_Sample/crr
      -- CP-element group 5: 	 call_stmt_261/call_stmt_261_Sample/$entry
      -- CP-element group 5: 	 call_stmt_261/call_stmt_261_sample_start_
      -- 
    crr_507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule_maxPool_CP_488_elements(5), ack => call_stmt_261_call_req_0); -- 
    readModule_maxPool_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "readModule_maxPool_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule_maxPool_CP_488_elements(1) & readModule_maxPool_CP_488_elements(7);
      gj_readModule_maxPool_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule_maxPool_CP_488_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	8 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 call_stmt_261/call_stmt_261_Update/ccr
      -- CP-element group 6: 	 call_stmt_261/call_stmt_261_Update/$entry
      -- CP-element group 6: 	 call_stmt_261/call_stmt_261_update_start_
      -- 
    ccr_512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule_maxPool_CP_488_elements(6), ack => call_stmt_261_call_req_1); -- 
    readModule_maxPool_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "readModule_maxPool_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule_maxPool_CP_488_elements(4) & readModule_maxPool_CP_488_elements(8);
      gj_readModule_maxPool_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule_maxPool_CP_488_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: successors 
    -- CP-element group 7: marked-successors 
    -- CP-element group 7: 	3 
    -- CP-element group 7: 	5 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_261/call_stmt_261_Sample/cra
      -- CP-element group 7: 	 call_stmt_261/call_stmt_261_Sample/$exit
      -- CP-element group 7: 	 call_stmt_261/call_stmt_261_sample_completed_
      -- 
    cra_508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_261_call_ack_0, ack => readModule_maxPool_CP_488_elements(7)); -- 
    -- CP-element group 8:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	12 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	6 
    -- CP-element group 8:  members (4) 
      -- CP-element group 8: 	 call_stmt_261/$exit
      -- CP-element group 8: 	 call_stmt_261/call_stmt_261_Update/cca
      -- CP-element group 8: 	 call_stmt_261/call_stmt_261_Update/$exit
      -- CP-element group 8: 	 call_stmt_261/call_stmt_261_update_completed_
      -- 
    cca_513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_261_call_ack_1, ack => readModule_maxPool_CP_488_elements(8)); -- 
    -- CP-element group 9:  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 index_update_enable
      -- 
    readModule_maxPool_CP_488_elements(9) <= readModule_maxPool_CP_488_elements(2);
    -- CP-element group 10:  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	3 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 address_update_enable
      -- 
    readModule_maxPool_CP_488_elements(10) <= readModule_maxPool_CP_488_elements(3);
    -- CP-element group 11:  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	4 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 data_update_enable
      -- 
    -- CP-element group 12:  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	8 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 $exit
      -- 
    readModule_maxPool_CP_488_elements(12) <= readModule_maxPool_CP_488_elements(8);
    --  hookup: inputs to control-path 
    readModule_maxPool_CP_488_elements(11) <= data_update_enable;
    -- hookup: output from control-path 
    address_update_enable <= readModule_maxPool_CP_488_elements(10);
    index_update_enable <= readModule_maxPool_CP_488_elements(9);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_258_wire : std_logic_vector(31 downto 0);
    signal konst_255_wire_constant : std_logic_vector(0 downto 0);
    signal konst_256_wire_constant : std_logic_vector(31 downto 0);
    signal konst_259_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_255_wire_constant <= "1";
    konst_256_wire_constant <= "00000000000000000000000000000000";
    konst_259_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- binary operator ADD_u32_u32_258_inst
    process(address_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address_buffer, konst_256_wire_constant, tmp_var);
      ADD_u32_u32_258_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_261_call 
    memoryModule_call_group_0: Block -- 
      signal data_in: std_logic_vector(96 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_261_call_req_0;
      call_stmt_261_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_261_call_req_1;
      call_stmt_261_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      memoryModule_call_group_0_gI: SplitGuardInterface generic map(name => "memoryModule_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_255_wire_constant & ADD_u32_u32_258_wire & konst_259_wire_constant;
      data_buffer <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 97,
        owidth => 97,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => memoryModule_call_reqs(0),
          ackR => memoryModule_call_acks(0),
          dataR => memoryModule_call_data(96 downto 0),
          tagR => memoryModule_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => memoryModule_return_acks(0), -- cross-over
          ackL => memoryModule_return_reqs(0), -- cross-over
          dataL => memoryModule_return_data(63 downto 0),
          tagL => memoryModule_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end readModule_maxPool_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendOutput is -- 
  generic (tag_length : integer); 
  port ( -- 
    system_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    system_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    system_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    readModule1_call_reqs : out  std_logic_vector(0 downto 0);
    readModule1_call_acks : in   std_logic_vector(0 downto 0);
    readModule1_call_data : out  std_logic_vector(31 downto 0);
    readModule1_call_tag  :  out  std_logic_vector(0 downto 0);
    readModule1_return_reqs : out  std_logic_vector(0 downto 0);
    readModule1_return_acks : in   std_logic_vector(0 downto 0);
    readModule1_return_data : in   std_logic_vector(63 downto 0);
    readModule1_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendOutput;
architecture sendOutput_arch of sendOutput is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal sendOutput_CP_1671_start: Boolean;
  signal sendOutput_CP_1671_symbol: Boolean;
  -- volatile/operator module components. 
  component readModule1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      address : in  std_logic_vector(31 downto 0);
      data : out  std_logic_vector(63 downto 0);
      memoryModule_call_reqs : out  std_logic_vector(0 downto 0);
      memoryModule_call_acks : in   std_logic_vector(0 downto 0);
      memoryModule_call_data : out  std_logic_vector(96 downto 0);
      memoryModule_call_tag  :  out  std_logic_vector(0 downto 0);
      memoryModule_return_reqs : out  std_logic_vector(0 downto 0);
      memoryModule_return_acks : in   std_logic_vector(0 downto 0);
      memoryModule_return_data : in   std_logic_vector(63 downto 0);
      memoryModule_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal WPIPE_system_output_pipe_1133_inst_ack_0 : boolean;
  signal type_cast_1101_inst_ack_0 : boolean;
  signal WPIPE_system_output_pipe_1139_inst_req_0 : boolean;
  signal type_cast_1091_inst_req_1 : boolean;
  signal type_cast_1091_inst_req_0 : boolean;
  signal type_cast_1101_inst_req_0 : boolean;
  signal WPIPE_system_output_pipe_1136_inst_ack_1 : boolean;
  signal type_cast_1091_inst_ack_1 : boolean;
  signal type_cast_1131_inst_req_0 : boolean;
  signal WPIPE_system_output_pipe_1139_inst_ack_0 : boolean;
  signal WPIPE_system_output_pipe_1142_inst_req_1 : boolean;
  signal WPIPE_system_output_pipe_1151_inst_ack_0 : boolean;
  signal WPIPE_system_output_pipe_1142_inst_req_0 : boolean;
  signal call_stmt_1058_call_req_0 : boolean;
  signal type_cast_1061_inst_req_1 : boolean;
  signal type_cast_1111_inst_ack_1 : boolean;
  signal type_cast_1081_inst_ack_1 : boolean;
  signal WPIPE_system_output_pipe_1142_inst_ack_0 : boolean;
  signal type_cast_1061_inst_ack_1 : boolean;
  signal type_cast_1091_inst_ack_0 : boolean;
  signal type_cast_1111_inst_req_1 : boolean;
  signal type_cast_1081_inst_req_1 : boolean;
  signal WPIPE_system_output_pipe_1136_inst_req_1 : boolean;
  signal WPIPE_system_output_pipe_1139_inst_ack_1 : boolean;
  signal WPIPE_system_output_pipe_1151_inst_req_1 : boolean;
  signal type_cast_1061_inst_req_0 : boolean;
  signal type_cast_1061_inst_ack_0 : boolean;
  signal WPIPE_system_output_pipe_1148_inst_ack_1 : boolean;
  signal WPIPE_system_output_pipe_1133_inst_req_1 : boolean;
  signal WPIPE_system_output_pipe_1133_inst_req_0 : boolean;
  signal WPIPE_system_output_pipe_1139_inst_req_1 : boolean;
  signal WPIPE_system_output_pipe_1136_inst_ack_0 : boolean;
  signal type_cast_1111_inst_ack_0 : boolean;
  signal phi_stmt_1048_req_0 : boolean;
  signal WPIPE_system_output_pipe_1136_inst_req_0 : boolean;
  signal type_cast_1111_inst_req_0 : boolean;
  signal type_cast_1121_inst_ack_1 : boolean;
  signal type_cast_1081_inst_ack_0 : boolean;
  signal type_cast_1121_inst_req_1 : boolean;
  signal WPIPE_system_output_pipe_1145_inst_ack_1 : boolean;
  signal WPIPE_system_output_pipe_1148_inst_ack_0 : boolean;
  signal WPIPE_system_output_pipe_1145_inst_req_1 : boolean;
  signal WPIPE_system_output_pipe_1151_inst_req_0 : boolean;
  signal type_cast_1131_inst_ack_1 : boolean;
  signal WPIPE_system_output_pipe_1148_inst_req_0 : boolean;
  signal if_stmt_1169_branch_ack_1 : boolean;
  signal type_cast_1081_inst_req_0 : boolean;
  signal WPIPE_system_output_pipe_1148_inst_req_1 : boolean;
  signal if_stmt_1169_branch_ack_0 : boolean;
  signal type_cast_1131_inst_req_1 : boolean;
  signal type_cast_1121_inst_ack_0 : boolean;
  signal type_cast_1121_inst_req_0 : boolean;
  signal WPIPE_system_output_pipe_1145_inst_ack_0 : boolean;
  signal WPIPE_system_output_pipe_1145_inst_req_0 : boolean;
  signal call_stmt_1058_call_ack_1 : boolean;
  signal WPIPE_system_output_pipe_1142_inst_ack_1 : boolean;
  signal call_stmt_1058_call_req_1 : boolean;
  signal type_cast_1131_inst_ack_0 : boolean;
  signal phi_stmt_1048_req_1 : boolean;
  signal if_stmt_1169_branch_req_0 : boolean;
  signal call_stmt_1058_call_ack_0 : boolean;
  signal WPIPE_system_output_pipe_1151_inst_ack_1 : boolean;
  signal type_cast_1071_inst_ack_1 : boolean;
  signal WPIPE_system_output_pipe_1154_inst_ack_1 : boolean;
  signal WPIPE_system_output_pipe_1154_inst_req_1 : boolean;
  signal type_cast_1101_inst_ack_1 : boolean;
  signal type_cast_1101_inst_req_1 : boolean;
  signal type_cast_1071_inst_req_1 : boolean;
  signal WPIPE_system_output_pipe_1154_inst_ack_0 : boolean;
  signal phi_stmt_1048_ack_0 : boolean;
  signal type_cast_1054_inst_req_1 : boolean;
  signal type_cast_1054_inst_req_0 : boolean;
  signal type_cast_1054_inst_ack_0 : boolean;
  signal type_cast_1054_inst_ack_1 : boolean;
  signal WPIPE_system_output_pipe_1154_inst_req_0 : boolean;
  signal type_cast_1071_inst_ack_0 : boolean;
  signal type_cast_1071_inst_req_0 : boolean;
  signal WPIPE_system_output_pipe_1133_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendOutput_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendOutput_CP_1671_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendOutput_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_1671_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendOutput_CP_1671_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_1671_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendOutput_CP_1671: Block -- control-path 
    signal sendOutput_CP_1671_elements: BooleanArray(49 downto 0);
    -- 
  begin -- 
    sendOutput_CP_1671_elements(0) <= sendOutput_CP_1671_start;
    sendOutput_CP_1671_symbol <= sendOutput_CP_1671_elements(42);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	44 
    -- CP-element group 0:  members (7) 
      -- CP-element group 0: 	 branch_block_stmt_1045/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1045/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_1045/bbx_xnph_forx_xbody
      -- CP-element group 0: 	 branch_block_stmt_1045/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1048/phi_stmt_1048_sources/$entry
      -- CP-element group 0: 	 branch_block_stmt_1045/branch_block_stmt_1045__entry__
      -- CP-element group 0: 	 branch_block_stmt_1045/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1048/$entry
      -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	49 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/call_stmt_1058_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/call_stmt_1058_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/call_stmt_1058_Sample/cra
      -- 
    cra_1700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1058_call_ack_0, ack => sendOutput_CP_1671_elements(1)); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	49 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	17 
    -- CP-element group 2:  members (27) 
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1091_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1121_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1101_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1091_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1101_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1131_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1091_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/call_stmt_1058_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1071_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1101_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1131_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1061_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1061_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1131_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1111_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1081_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1111_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1121_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1081_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1061_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/call_stmt_1058_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1121_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1111_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1081_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/call_stmt_1058_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1071_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1071_Sample/$entry
      -- 
    cca_1705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1058_call_ack_1, ack => sendOutput_CP_1671_elements(2)); -- 
    rr_1713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(2), ack => type_cast_1061_inst_req_0); -- 
    rr_1727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(2), ack => type_cast_1071_inst_req_0); -- 
    rr_1741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(2), ack => type_cast_1081_inst_req_0); -- 
    rr_1755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(2), ack => type_cast_1091_inst_req_0); -- 
    rr_1769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(2), ack => type_cast_1101_inst_req_0); -- 
    rr_1783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(2), ack => type_cast_1111_inst_req_0); -- 
    rr_1797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(2), ack => type_cast_1121_inst_req_0); -- 
    rr_1811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(2), ack => type_cast_1131_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1061_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1061_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1061_sample_completed_
      -- 
    ra_1714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1061_inst_ack_0, ack => sendOutput_CP_1671_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	49 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	39 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1061_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1061_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1061_update_completed_
      -- 
    ca_1719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1061_inst_ack_1, ack => sendOutput_CP_1671_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1071_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1071_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1071_Sample/$exit
      -- 
    ra_1728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1071_inst_ack_0, ack => sendOutput_CP_1671_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	49 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	36 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1071_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1071_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1071_update_completed_
      -- 
    ca_1733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1071_inst_ack_1, ack => sendOutput_CP_1671_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1081_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1081_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1081_sample_completed_
      -- 
    ra_1742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1081_inst_ack_0, ack => sendOutput_CP_1671_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	49 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	33 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1081_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1081_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1081_update_completed_
      -- 
    ca_1747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1081_inst_ack_1, ack => sendOutput_CP_1671_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1091_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1091_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1091_Sample/ra
      -- 
    ra_1756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1091_inst_ack_0, ack => sendOutput_CP_1671_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	49 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	30 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1091_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1091_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1091_update_completed_
      -- 
    ca_1761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1091_inst_ack_1, ack => sendOutput_CP_1671_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1101_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1101_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1101_sample_completed_
      -- 
    ra_1770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1101_inst_ack_0, ack => sendOutput_CP_1671_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	49 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	27 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1101_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1101_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1101_Update/$exit
      -- 
    ca_1775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1101_inst_ack_1, ack => sendOutput_CP_1671_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1111_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1111_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1111_sample_completed_
      -- 
    ra_1784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1111_inst_ack_0, ack => sendOutput_CP_1671_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	49 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	24 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1111_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1111_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1111_update_completed_
      -- 
    ca_1789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1111_inst_ack_1, ack => sendOutput_CP_1671_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1121_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1121_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1121_Sample/$exit
      -- 
    ra_1798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1121_inst_ack_0, ack => sendOutput_CP_1671_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	49 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	21 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1121_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1121_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1121_update_completed_
      -- 
    ca_1803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1121_inst_ack_1, ack => sendOutput_CP_1671_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1131_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1131_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1131_Sample/ra
      -- 
    ra_1812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1131_inst_ack_0, ack => sendOutput_CP_1671_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	49 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1131_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1133_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1133_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1133_Sample/req
      -- CP-element group 18: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1131_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1131_Update/$exit
      -- 
    ca_1817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1131_inst_ack_1, ack => sendOutput_CP_1671_elements(18)); -- 
    req_1825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(18), ack => WPIPE_system_output_pipe_1133_inst_req_0); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1133_Sample/ack
      -- CP-element group 19: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1133_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1133_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1133_Update/req
      -- CP-element group 19: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1133_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1133_update_start_
      -- 
    ack_1826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1133_inst_ack_0, ack => sendOutput_CP_1671_elements(19)); -- 
    req_1830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(19), ack => WPIPE_system_output_pipe_1133_inst_req_1); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1133_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1133_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1133_Update/ack
      -- 
    ack_1831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1133_inst_ack_1, ack => sendOutput_CP_1671_elements(20)); -- 
    -- CP-element group 21:  join  transition  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	16 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1136_Sample/req
      -- CP-element group 21: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1136_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1136_sample_start_
      -- 
    req_1839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(21), ack => WPIPE_system_output_pipe_1136_inst_req_0); -- 
    sendOutput_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_1671_elements(16) & sendOutput_CP_1671_elements(20);
      gj_sendOutput_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_1671_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1136_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1136_Update/req
      -- CP-element group 22: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1136_Sample/ack
      -- CP-element group 22: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1136_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1136_update_start_
      -- CP-element group 22: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1136_sample_completed_
      -- 
    ack_1840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1136_inst_ack_0, ack => sendOutput_CP_1671_elements(22)); -- 
    req_1844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(22), ack => WPIPE_system_output_pipe_1136_inst_req_1); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1136_Update/ack
      -- CP-element group 23: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1136_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1136_update_completed_
      -- 
    ack_1845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1136_inst_ack_1, ack => sendOutput_CP_1671_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	14 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1139_Sample/req
      -- CP-element group 24: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1139_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1139_sample_start_
      -- 
    req_1853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(24), ack => WPIPE_system_output_pipe_1139_inst_req_0); -- 
    sendOutput_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_1671_elements(14) & sendOutput_CP_1671_elements(23);
      gj_sendOutput_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_1671_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1139_Sample/ack
      -- CP-element group 25: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1139_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1139_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1139_Update/req
      -- CP-element group 25: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1139_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1139_sample_completed_
      -- 
    ack_1854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1139_inst_ack_0, ack => sendOutput_CP_1671_elements(25)); -- 
    req_1858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(25), ack => WPIPE_system_output_pipe_1139_inst_req_1); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1139_Update/ack
      -- CP-element group 26: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1139_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1139_update_completed_
      -- 
    ack_1859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1139_inst_ack_1, ack => sendOutput_CP_1671_elements(26)); -- 
    -- CP-element group 27:  join  transition  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	12 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1142_Sample/req
      -- CP-element group 27: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1142_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1142_sample_start_
      -- 
    req_1867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(27), ack => WPIPE_system_output_pipe_1142_inst_req_0); -- 
    sendOutput_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_1671_elements(12) & sendOutput_CP_1671_elements(26);
      gj_sendOutput_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_1671_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1142_Update/req
      -- CP-element group 28: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1142_Sample/ack
      -- CP-element group 28: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1142_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1142_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1142_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1142_Update/$entry
      -- 
    ack_1868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1142_inst_ack_0, ack => sendOutput_CP_1671_elements(28)); -- 
    req_1872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(28), ack => WPIPE_system_output_pipe_1142_inst_req_1); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1142_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1142_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1142_Update/ack
      -- 
    ack_1873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1142_inst_ack_1, ack => sendOutput_CP_1671_elements(29)); -- 
    -- CP-element group 30:  join  transition  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	10 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1145_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1145_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1145_Sample/req
      -- 
    req_1881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(30), ack => WPIPE_system_output_pipe_1145_inst_req_0); -- 
    sendOutput_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_1671_elements(10) & sendOutput_CP_1671_elements(29);
      gj_sendOutput_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_1671_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1145_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1145_update_start_
      -- CP-element group 31: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1145_Update/req
      -- CP-element group 31: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1145_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1145_Sample/ack
      -- CP-element group 31: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1145_Sample/$exit
      -- 
    ack_1882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1145_inst_ack_0, ack => sendOutput_CP_1671_elements(31)); -- 
    req_1886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(31), ack => WPIPE_system_output_pipe_1145_inst_req_1); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1145_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1145_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1145_Update/ack
      -- 
    ack_1887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1145_inst_ack_1, ack => sendOutput_CP_1671_elements(32)); -- 
    -- CP-element group 33:  join  transition  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	8 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1148_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1148_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1148_Sample/req
      -- 
    req_1895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(33), ack => WPIPE_system_output_pipe_1148_inst_req_0); -- 
    sendOutput_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_1671_elements(8) & sendOutput_CP_1671_elements(32);
      gj_sendOutput_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_1671_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1148_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1148_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1148_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1148_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1148_Sample/ack
      -- CP-element group 34: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1148_Update/req
      -- 
    ack_1896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1148_inst_ack_0, ack => sendOutput_CP_1671_elements(34)); -- 
    req_1900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(34), ack => WPIPE_system_output_pipe_1148_inst_req_1); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1148_Update/ack
      -- CP-element group 35: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1148_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1148_update_completed_
      -- 
    ack_1901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1148_inst_ack_1, ack => sendOutput_CP_1671_elements(35)); -- 
    -- CP-element group 36:  join  transition  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	6 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1151_Sample/req
      -- CP-element group 36: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1151_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1151_sample_start_
      -- 
    req_1909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(36), ack => WPIPE_system_output_pipe_1151_inst_req_0); -- 
    sendOutput_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_1671_elements(6) & sendOutput_CP_1671_elements(35);
      gj_sendOutput_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_1671_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1151_Sample/ack
      -- CP-element group 37: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1151_Update/req
      -- CP-element group 37: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1151_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1151_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1151_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1151_update_start_
      -- 
    ack_1910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1151_inst_ack_0, ack => sendOutput_CP_1671_elements(37)); -- 
    req_1914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(37), ack => WPIPE_system_output_pipe_1151_inst_req_1); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1151_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1151_Update/ack
      -- CP-element group 38: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1151_update_completed_
      -- 
    ack_1915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1151_inst_ack_1, ack => sendOutput_CP_1671_elements(38)); -- 
    -- CP-element group 39:  join  transition  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	4 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1154_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1154_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1154_Sample/req
      -- 
    req_1923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(39), ack => WPIPE_system_output_pipe_1154_inst_req_0); -- 
    sendOutput_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_1671_elements(4) & sendOutput_CP_1671_elements(38);
      gj_sendOutput_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_1671_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (6) 
      -- CP-element group 40: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1154_update_start_
      -- CP-element group 40: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1154_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1154_Update/req
      -- CP-element group 40: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1154_Update/$entry
      -- CP-element group 40: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1154_Sample/ack
      -- CP-element group 40: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1154_Sample/$exit
      -- 
    ack_1924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1154_inst_ack_0, ack => sendOutput_CP_1671_elements(40)); -- 
    req_1928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(40), ack => WPIPE_system_output_pipe_1154_inst_req_1); -- 
    -- CP-element group 41:  branch  transition  place  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (13) 
      -- CP-element group 41: 	 branch_block_stmt_1045/if_stmt_1169__entry__
      -- CP-element group 41: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168__exit__
      -- CP-element group 41: 	 branch_block_stmt_1045/if_stmt_1169_if_link/$entry
      -- CP-element group 41: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/$exit
      -- CP-element group 41: 	 branch_block_stmt_1045/R_exitcond1_1170_place
      -- CP-element group 41: 	 branch_block_stmt_1045/if_stmt_1169_eval_test/branch_req
      -- CP-element group 41: 	 branch_block_stmt_1045/if_stmt_1169_eval_test/$exit
      -- CP-element group 41: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1154_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1045/if_stmt_1169_eval_test/$entry
      -- CP-element group 41: 	 branch_block_stmt_1045/if_stmt_1169_dead_link/$entry
      -- CP-element group 41: 	 branch_block_stmt_1045/if_stmt_1169_else_link/$entry
      -- CP-element group 41: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1154_Update/ack
      -- CP-element group 41: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/WPIPE_system_output_pipe_1154_Update/$exit
      -- 
    ack_1929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1154_inst_ack_1, ack => sendOutput_CP_1671_elements(41)); -- 
    branch_req_1937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(41), ack => if_stmt_1169_branch_req_0); -- 
    -- CP-element group 42:  merge  transition  place  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (21) 
      -- CP-element group 42: 	 $exit
      -- CP-element group 42: 	 branch_block_stmt_1045/if_stmt_1169_if_link/$exit
      -- CP-element group 42: 	 branch_block_stmt_1045/forx_xbody_forx_xend_PhiReq/$exit
      -- CP-element group 42: 	 branch_block_stmt_1045/merge_stmt_1175_PhiReqMerge
      -- CP-element group 42: 	 branch_block_stmt_1045/merge_stmt_1175_PhiAck/$entry
      -- CP-element group 42: 	 branch_block_stmt_1045/merge_stmt_1175_PhiAck/$exit
      -- CP-element group 42: 	 branch_block_stmt_1045/merge_stmt_1175_PhiAck/dummy
      -- CP-element group 42: 	 branch_block_stmt_1045/branch_block_stmt_1045__exit__
      -- CP-element group 42: 	 branch_block_stmt_1045/merge_stmt_1177_PhiReqMerge
      -- CP-element group 42: 	 branch_block_stmt_1045/return___PhiReq/$entry
      -- CP-element group 42: 	 branch_block_stmt_1045/return___PhiReq/$exit
      -- CP-element group 42: 	 branch_block_stmt_1045/if_stmt_1169_if_link/if_choice_transition
      -- CP-element group 42: 	 branch_block_stmt_1045/merge_stmt_1177__exit__
      -- CP-element group 42: 	 branch_block_stmt_1045/return__
      -- CP-element group 42: 	 branch_block_stmt_1045/merge_stmt_1175__exit__
      -- CP-element group 42: 	 branch_block_stmt_1045/$exit
      -- CP-element group 42: 	 branch_block_stmt_1045/forx_xbody_forx_xend
      -- CP-element group 42: 	 branch_block_stmt_1045/forx_xbody_forx_xend_PhiReq/$entry
      -- CP-element group 42: 	 branch_block_stmt_1045/merge_stmt_1177_PhiAck/$entry
      -- CP-element group 42: 	 branch_block_stmt_1045/merge_stmt_1177_PhiAck/$exit
      -- CP-element group 42: 	 branch_block_stmt_1045/merge_stmt_1177_PhiAck/dummy
      -- 
    if_choice_transition_1942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1169_branch_ack_1, ack => sendOutput_CP_1671_elements(42)); -- 
    -- CP-element group 43:  fork  transition  place  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43: 	46 
    -- CP-element group 43:  members (12) 
      -- CP-element group 43: 	 branch_block_stmt_1045/forx_xbody_forx_xbody_PhiReq/phi_stmt_1048/$entry
      -- CP-element group 43: 	 branch_block_stmt_1045/forx_xbody_forx_xbody_PhiReq/phi_stmt_1048/phi_stmt_1048_sources/type_cast_1054/$entry
      -- CP-element group 43: 	 branch_block_stmt_1045/forx_xbody_forx_xbody_PhiReq/phi_stmt_1048/phi_stmt_1048_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1045/if_stmt_1169_else_link/else_choice_transition
      -- CP-element group 43: 	 branch_block_stmt_1045/forx_xbody_forx_xbody_PhiReq/phi_stmt_1048/phi_stmt_1048_sources/type_cast_1054/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_1045/forx_xbody_forx_xbody_PhiReq/phi_stmt_1048/phi_stmt_1048_sources/type_cast_1054/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1045/forx_xbody_forx_xbody
      -- CP-element group 43: 	 branch_block_stmt_1045/if_stmt_1169_else_link/$exit
      -- CP-element group 43: 	 branch_block_stmt_1045/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1045/forx_xbody_forx_xbody_PhiReq/phi_stmt_1048/phi_stmt_1048_sources/type_cast_1054/SplitProtocol/Update/cr
      -- CP-element group 43: 	 branch_block_stmt_1045/forx_xbody_forx_xbody_PhiReq/phi_stmt_1048/phi_stmt_1048_sources/type_cast_1054/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1045/forx_xbody_forx_xbody_PhiReq/phi_stmt_1048/phi_stmt_1048_sources/type_cast_1054/SplitProtocol/Sample/rr
      -- 
    else_choice_transition_1946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1169_branch_ack_0, ack => sendOutput_CP_1671_elements(43)); -- 
    cr_1983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(43), ack => type_cast_1054_inst_req_1); -- 
    rr_1978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(43), ack => type_cast_1054_inst_req_0); -- 
    -- CP-element group 44:  transition  output  delay-element  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	48 
    -- CP-element group 44:  members (5) 
      -- CP-element group 44: 	 branch_block_stmt_1045/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1048/phi_stmt_1048_req
      -- CP-element group 44: 	 branch_block_stmt_1045/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1048/phi_stmt_1048_sources/type_cast_1052_konst_delay_trans
      -- CP-element group 44: 	 branch_block_stmt_1045/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1048/phi_stmt_1048_sources/$exit
      -- CP-element group 44: 	 branch_block_stmt_1045/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1048/$exit
      -- CP-element group 44: 	 branch_block_stmt_1045/bbx_xnph_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_1048_req_1959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1048_req_1959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(44), ack => phi_stmt_1048_req_0); -- 
    -- Element group sendOutput_CP_1671_elements(44) is a control-delay.
    cp_element_44_delay: control_delay_element  generic map(name => " 44_delay", delay_value => 1)  port map(req => sendOutput_CP_1671_elements(0), ack => sendOutput_CP_1671_elements(44), clk => clk, reset =>reset);
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_1045/forx_xbody_forx_xbody_PhiReq/phi_stmt_1048/phi_stmt_1048_sources/type_cast_1054/SplitProtocol/Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1045/forx_xbody_forx_xbody_PhiReq/phi_stmt_1048/phi_stmt_1048_sources/type_cast_1054/SplitProtocol/Sample/ra
      -- 
    ra_1979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1054_inst_ack_0, ack => sendOutput_CP_1671_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	43 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1045/forx_xbody_forx_xbody_PhiReq/phi_stmt_1048/phi_stmt_1048_sources/type_cast_1054/SplitProtocol/Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1045/forx_xbody_forx_xbody_PhiReq/phi_stmt_1048/phi_stmt_1048_sources/type_cast_1054/SplitProtocol/Update/ca
      -- 
    ca_1984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1054_inst_ack_1, ack => sendOutput_CP_1671_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (6) 
      -- CP-element group 47: 	 branch_block_stmt_1045/forx_xbody_forx_xbody_PhiReq/phi_stmt_1048/$exit
      -- CP-element group 47: 	 branch_block_stmt_1045/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 47: 	 branch_block_stmt_1045/forx_xbody_forx_xbody_PhiReq/phi_stmt_1048/phi_stmt_1048_sources/type_cast_1054/SplitProtocol/$exit
      -- CP-element group 47: 	 branch_block_stmt_1045/forx_xbody_forx_xbody_PhiReq/phi_stmt_1048/phi_stmt_1048_req
      -- CP-element group 47: 	 branch_block_stmt_1045/forx_xbody_forx_xbody_PhiReq/phi_stmt_1048/phi_stmt_1048_sources/$exit
      -- CP-element group 47: 	 branch_block_stmt_1045/forx_xbody_forx_xbody_PhiReq/phi_stmt_1048/phi_stmt_1048_sources/type_cast_1054/$exit
      -- 
    phi_stmt_1048_req_1985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1048_req_1985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(47), ack => phi_stmt_1048_req_1); -- 
    sendOutput_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_1671_elements(45) & sendOutput_CP_1671_elements(46);
      gj_sendOutput_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_1671_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  merge  transition  place  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	44 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_1045/merge_stmt_1047_PhiReqMerge
      -- CP-element group 48: 	 branch_block_stmt_1045/merge_stmt_1047_PhiAck/$entry
      -- 
    sendOutput_CP_1671_elements(48) <= OrReduce(sendOutput_CP_1671_elements(44) & sendOutput_CP_1671_elements(47));
    -- CP-element group 49:  fork  transition  place  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	1 
    -- CP-element group 49: 	2 
    -- CP-element group 49: 	4 
    -- CP-element group 49: 	6 
    -- CP-element group 49: 	8 
    -- CP-element group 49: 	10 
    -- CP-element group 49: 	12 
    -- CP-element group 49: 	14 
    -- CP-element group 49: 	16 
    -- CP-element group 49: 	18 
    -- CP-element group 49:  members (35) 
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1091_Update/cr
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168__entry__
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1061_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1101_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/call_stmt_1058_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1071_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1121_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1045/merge_stmt_1047__exit__
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1111_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/call_stmt_1058_Sample/crr
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1061_Update/cr
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1091_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1091_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1111_Update/cr
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1101_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/call_stmt_1058_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1081_Update/cr
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1131_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/$entry
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/call_stmt_1058_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1081_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1121_Update/cr
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1131_Update/cr
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1061_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1111_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1121_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1081_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1131_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/call_stmt_1058_Update/ccr
      -- CP-element group 49: 	 branch_block_stmt_1045/merge_stmt_1047_PhiAck/$exit
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/call_stmt_1058_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1101_Update/cr
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1071_Update/cr
      -- CP-element group 49: 	 branch_block_stmt_1045/merge_stmt_1047_PhiAck/phi_stmt_1048_ack
      -- CP-element group 49: 	 branch_block_stmt_1045/call_stmt_1058_to_assign_stmt_1168/type_cast_1071_Update/$entry
      -- 
    phi_stmt_1048_ack_1990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1048_ack_0, ack => sendOutput_CP_1671_elements(49)); -- 
    cr_1760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(49), ack => type_cast_1091_inst_req_1); -- 
    crr_1699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(49), ack => call_stmt_1058_call_req_0); -- 
    cr_1718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(49), ack => type_cast_1061_inst_req_1); -- 
    cr_1788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(49), ack => type_cast_1111_inst_req_1); -- 
    cr_1746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(49), ack => type_cast_1081_inst_req_1); -- 
    cr_1802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(49), ack => type_cast_1121_inst_req_1); -- 
    cr_1816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(49), ack => type_cast_1131_inst_req_1); -- 
    ccr_1704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(49), ack => call_stmt_1058_call_req_1); -- 
    cr_1774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(49), ack => type_cast_1101_inst_req_1); -- 
    cr_1732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_1671_elements(49), ack => type_cast_1071_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal call_1058 : std_logic_vector(63 downto 0);
    signal conv14_1082 : std_logic_vector(7 downto 0);
    signal conv20_1092 : std_logic_vector(7 downto 0);
    signal conv26_1102 : std_logic_vector(7 downto 0);
    signal conv32_1112 : std_logic_vector(7 downto 0);
    signal conv38_1122 : std_logic_vector(7 downto 0);
    signal conv44_1132 : std_logic_vector(7 downto 0);
    signal conv8_1072 : std_logic_vector(7 downto 0);
    signal conv_1062 : std_logic_vector(7 downto 0);
    signal exitcond1_1168 : std_logic_vector(0 downto 0);
    signal iNsTr_1_1048 : std_logic_vector(31 downto 0);
    signal inc_1162 : std_logic_vector(31 downto 0);
    signal shr11_1078 : std_logic_vector(63 downto 0);
    signal shr17_1088 : std_logic_vector(63 downto 0);
    signal shr23_1098 : std_logic_vector(63 downto 0);
    signal shr29_1108 : std_logic_vector(63 downto 0);
    signal shr35_1118 : std_logic_vector(63 downto 0);
    signal shr41_1128 : std_logic_vector(63 downto 0);
    signal shr_1068 : std_logic_vector(63 downto 0);
    signal type_cast_1052_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1054_wire : std_logic_vector(31 downto 0);
    signal type_cast_1066_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1076_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1086_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1096_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1106_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1116_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1126_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1160_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1166_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    type_cast_1052_wire_constant <= "00000000000000000000000000000000";
    type_cast_1066_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1076_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1086_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1096_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1106_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1116_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1126_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1160_wire_constant <= "00000000000000000000000000000001";
    type_cast_1166_wire_constant <= "00000000000000001100010000000000";
    phi_stmt_1048: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1052_wire_constant & type_cast_1054_wire;
      req <= phi_stmt_1048_req_0 & phi_stmt_1048_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1048",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1048_ack_0,
          idata => idata,
          odata => iNsTr_1_1048,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1048
    type_cast_1054_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1054_inst_req_0;
      type_cast_1054_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1054_inst_req_1;
      type_cast_1054_inst_ack_1<= rack(0);
      type_cast_1054_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1054_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_1162,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1054_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1061_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1061_inst_req_0;
      type_cast_1061_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1061_inst_req_1;
      type_cast_1061_inst_ack_1<= rack(0);
      type_cast_1061_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1061_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1058,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1062,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1071_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1071_inst_req_0;
      type_cast_1071_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1071_inst_req_1;
      type_cast_1071_inst_ack_1<= rack(0);
      type_cast_1071_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1071_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_1068,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_1072,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1081_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1081_inst_req_0;
      type_cast_1081_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1081_inst_req_1;
      type_cast_1081_inst_ack_1<= rack(0);
      type_cast_1081_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1081_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr11_1078,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv14_1082,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1091_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1091_inst_req_0;
      type_cast_1091_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1091_inst_req_1;
      type_cast_1091_inst_ack_1<= rack(0);
      type_cast_1091_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1091_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr17_1088,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_1092,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1101_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1101_inst_req_0;
      type_cast_1101_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1101_inst_req_1;
      type_cast_1101_inst_ack_1<= rack(0);
      type_cast_1101_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1101_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr23_1098,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_1102,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1111_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1111_inst_req_0;
      type_cast_1111_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1111_inst_req_1;
      type_cast_1111_inst_ack_1<= rack(0);
      type_cast_1111_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1111_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr29_1108,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_1112,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1121_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1121_inst_req_0;
      type_cast_1121_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1121_inst_req_1;
      type_cast_1121_inst_ack_1<= rack(0);
      type_cast_1121_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1121_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr35_1118,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_1122,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1131_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1131_inst_req_0;
      type_cast_1131_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1131_inst_req_1;
      type_cast_1131_inst_ack_1<= rack(0);
      type_cast_1131_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1131_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr41_1128,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_1132,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    if_stmt_1169_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1168;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1169_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1169_branch_req_0,
          ack0 => if_stmt_1169_branch_ack_0,
          ack1 => if_stmt_1169_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1161_inst
    process(iNsTr_1_1048) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_1_1048, type_cast_1160_wire_constant, tmp_var);
      inc_1162 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1167_inst
    process(inc_1162) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_1162, type_cast_1166_wire_constant, tmp_var);
      exitcond1_1168 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1067_inst
    process(call_1058) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1058, type_cast_1066_wire_constant, tmp_var);
      shr_1068 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1077_inst
    process(call_1058) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1058, type_cast_1076_wire_constant, tmp_var);
      shr11_1078 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1087_inst
    process(call_1058) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1058, type_cast_1086_wire_constant, tmp_var);
      shr17_1088 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1097_inst
    process(call_1058) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1058, type_cast_1096_wire_constant, tmp_var);
      shr23_1098 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1107_inst
    process(call_1058) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1058, type_cast_1106_wire_constant, tmp_var);
      shr29_1108 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1117_inst
    process(call_1058) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1058, type_cast_1116_wire_constant, tmp_var);
      shr35_1118 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1127_inst
    process(call_1058) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1058, type_cast_1126_wire_constant, tmp_var);
      shr41_1128 <= tmp_var; --
    end process;
    -- shared outport operator group (0) : WPIPE_system_output_pipe_1133_inst WPIPE_system_output_pipe_1136_inst WPIPE_system_output_pipe_1139_inst WPIPE_system_output_pipe_1142_inst WPIPE_system_output_pipe_1145_inst WPIPE_system_output_pipe_1148_inst WPIPE_system_output_pipe_1151_inst WPIPE_system_output_pipe_1154_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_system_output_pipe_1133_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_system_output_pipe_1136_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_system_output_pipe_1139_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_system_output_pipe_1142_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_system_output_pipe_1145_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_system_output_pipe_1148_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_system_output_pipe_1151_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_system_output_pipe_1154_inst_req_0;
      WPIPE_system_output_pipe_1133_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_system_output_pipe_1136_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_system_output_pipe_1139_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_system_output_pipe_1142_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_system_output_pipe_1145_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_system_output_pipe_1148_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_system_output_pipe_1151_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_system_output_pipe_1154_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_system_output_pipe_1133_inst_req_1;
      update_req_unguarded(6) <= WPIPE_system_output_pipe_1136_inst_req_1;
      update_req_unguarded(5) <= WPIPE_system_output_pipe_1139_inst_req_1;
      update_req_unguarded(4) <= WPIPE_system_output_pipe_1142_inst_req_1;
      update_req_unguarded(3) <= WPIPE_system_output_pipe_1145_inst_req_1;
      update_req_unguarded(2) <= WPIPE_system_output_pipe_1148_inst_req_1;
      update_req_unguarded(1) <= WPIPE_system_output_pipe_1151_inst_req_1;
      update_req_unguarded(0) <= WPIPE_system_output_pipe_1154_inst_req_1;
      WPIPE_system_output_pipe_1133_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_system_output_pipe_1136_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_system_output_pipe_1139_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_system_output_pipe_1142_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_system_output_pipe_1145_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_system_output_pipe_1148_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_system_output_pipe_1151_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_system_output_pipe_1154_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv44_1132 & conv38_1122 & conv32_1112 & conv26_1102 & conv20_1092 & conv14_1082 & conv8_1072 & conv_1062;
      system_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "system_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      system_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "system_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => system_output_pipe_pipe_write_req(0),
          oack => system_output_pipe_pipe_write_ack(0),
          odata => system_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1058_call 
    readModule1_call_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1058_call_req_0;
      call_stmt_1058_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1058_call_req_1;
      call_stmt_1058_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      readModule1_call_group_0_gI: SplitGuardInterface generic map(name => "readModule1_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= iNsTr_1_1048;
      call_1058 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 32,
        owidth => 32,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => readModule1_call_reqs(0),
          ackR => readModule1_call_acks(0),
          dataR => readModule1_call_data(31 downto 0),
          tagR => readModule1_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => readModule1_return_acks(0), -- cross-over
          ackL => readModule1_return_reqs(0), -- cross-over
          dataL => readModule1_return_data(63 downto 0),
          tagL => readModule1_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end sendOutput_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity systemTOP is -- 
  generic (tag_length : integer); 
  port ( -- 
    system_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    system_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    system_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    fill_input_call_reqs : out  std_logic_vector(0 downto 0);
    fill_input_call_acks : in   std_logic_vector(0 downto 0);
    fill_input_call_tag  :  out  std_logic_vector(0 downto 0);
    fill_input_return_reqs : out  std_logic_vector(0 downto 0);
    fill_input_return_acks : in   std_logic_vector(0 downto 0);
    fill_input_return_tag :  in   std_logic_vector(0 downto 0);
    maxPool4_call_reqs : out  std_logic_vector(0 downto 0);
    maxPool4_call_acks : in   std_logic_vector(0 downto 0);
    maxPool4_call_data : out  std_logic_vector(175 downto 0);
    maxPool4_call_tag  :  out  std_logic_vector(0 downto 0);
    maxPool4_return_reqs : out  std_logic_vector(0 downto 0);
    maxPool4_return_acks : in   std_logic_vector(0 downto 0);
    maxPool4_return_data : in   std_logic_vector(7 downto 0);
    maxPool4_return_tag :  in   std_logic_vector(0 downto 0);
    sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_call_acks : in   std_logic_vector(0 downto 0);
    sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
    sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_return_acks : in   std_logic_vector(0 downto 0);
    sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity systemTOP;
architecture systemTOP_arch of systemTOP is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal systemTOP_CP_2045_start: Boolean;
  signal systemTOP_CP_2045_symbol: Boolean;
  -- volatile/operator module components. 
  component fill_input is -- 
    generic (tag_length : integer); 
    port ( -- 
      system_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      system_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      system_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      writeModule1_call_reqs : out  std_logic_vector(0 downto 0);
      writeModule1_call_acks : in   std_logic_vector(0 downto 0);
      writeModule1_call_data : out  std_logic_vector(95 downto 0);
      writeModule1_call_tag  :  out  std_logic_vector(0 downto 0);
      writeModule1_return_reqs : out  std_logic_vector(0 downto 0);
      writeModule1_return_acks : in   std_logic_vector(0 downto 0);
      writeModule1_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component maxPool4 is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(31 downto 0);
      addr1 : in  std_logic_vector(31 downto 0);
      addr2 : in  std_logic_vector(31 downto 0);
      addr3 : in  std_logic_vector(31 downto 0);
      addr4 : in  std_logic_vector(31 downto 0);
      index1 : in  std_logic_vector(7 downto 0);
      index2 : in  std_logic_vector(7 downto 0);
      output : out  std_logic_vector(7 downto 0);
      readModule_maxPool_call_reqs : out  std_logic_vector(0 downto 0);
      readModule_maxPool_call_acks : in   std_logic_vector(0 downto 0);
      readModule_maxPool_call_data : out  std_logic_vector(39 downto 0);
      readModule_maxPool_call_tag  :  out  std_logic_vector(2 downto 0);
      readModule_maxPool_return_reqs : out  std_logic_vector(0 downto 0);
      readModule_maxPool_return_acks : in   std_logic_vector(0 downto 0);
      readModule_maxPool_return_data : in   std_logic_vector(63 downto 0);
      readModule_maxPool_return_tag :  in   std_logic_vector(2 downto 0);
      writeModule_maxPool_call_reqs : out  std_logic_vector(0 downto 0);
      writeModule_maxPool_call_acks : in   std_logic_vector(0 downto 0);
      writeModule_maxPool_call_data : out  std_logic_vector(103 downto 0);
      writeModule_maxPool_call_tag  :  out  std_logic_vector(0 downto 0);
      writeModule_maxPool_return_reqs : out  std_logic_vector(0 downto 0);
      writeModule_maxPool_return_acks : in   std_logic_vector(0 downto 0);
      writeModule_maxPool_return_data : in   std_logic_vector(0 downto 0);
      writeModule_maxPool_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      system_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      system_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      system_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      readModule1_call_reqs : out  std_logic_vector(0 downto 0);
      readModule1_call_acks : in   std_logic_vector(0 downto 0);
      readModule1_call_data : out  std_logic_vector(31 downto 0);
      readModule1_call_tag  :  out  std_logic_vector(0 downto 0);
      readModule1_return_reqs : out  std_logic_vector(0 downto 0);
      readModule1_return_acks : in   std_logic_vector(0 downto 0);
      readModule1_return_data : in   std_logic_vector(63 downto 0);
      readModule1_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal type_cast_1243_inst_req_1 : boolean;
  signal type_cast_1243_inst_ack_1 : boolean;
  signal type_cast_1233_inst_req_1 : boolean;
  signal W_colx_x1x_xi_1307_delayed_1_0_1323_inst_ack_1 : boolean;
  signal type_cast_1247_inst_req_1 : boolean;
  signal type_cast_1233_inst_ack_1 : boolean;
  signal type_cast_1238_inst_req_0 : boolean;
  signal type_cast_1247_inst_ack_1 : boolean;
  signal type_cast_1321_inst_req_1 : boolean;
  signal phi_stmt_1235_req_0 : boolean;
  signal type_cast_1321_inst_ack_1 : boolean;
  signal W_row18x_x1x_xi_1329_delayed_2_0_1348_inst_ack_1 : boolean;
  signal type_cast_1243_inst_req_0 : boolean;
  signal type_cast_1251_inst_req_1 : boolean;
  signal W_iNsTr_2_1278_delayed_1_0_1293_inst_req_1 : boolean;
  signal type_cast_1233_inst_req_0 : boolean;
  signal W_colx_x1x_xi_1307_delayed_1_0_1323_inst_req_1 : boolean;
  signal type_cast_1238_inst_ack_0 : boolean;
  signal type_cast_1247_inst_ack_0 : boolean;
  signal type_cast_1251_inst_ack_1 : boolean;
  signal type_cast_1228_inst_req_1 : boolean;
  signal type_cast_1247_inst_req_0 : boolean;
  signal type_cast_1251_inst_ack_0 : boolean;
  signal type_cast_1321_inst_req_0 : boolean;
  signal phi_stmt_1235_ack_0 : boolean;
  signal type_cast_1233_inst_ack_0 : boolean;
  signal phi_stmt_1235_req_1 : boolean;
  signal W_iNsTr_2_1278_delayed_1_0_1293_inst_ack_1 : boolean;
  signal W_colx_x1x_xi_1307_delayed_1_0_1323_inst_ack_0 : boolean;
  signal W_colx_x1x_xi_1307_delayed_1_0_1323_inst_req_0 : boolean;
  signal phi_stmt_1230_ack_0 : boolean;
  signal type_cast_1243_inst_ack_0 : boolean;
  signal type_cast_1321_inst_ack_0 : boolean;
  signal type_cast_1228_inst_ack_1 : boolean;
  signal W_iNsTr_2_1278_delayed_1_0_1293_inst_req_0 : boolean;
  signal type_cast_1346_inst_req_1 : boolean;
  signal W_row18x_x1x_xi_1329_delayed_2_0_1348_inst_req_1 : boolean;
  signal type_cast_1395_inst_ack_0 : boolean;
  signal type_cast_1399_inst_req_0 : boolean;
  signal type_cast_1399_inst_ack_0 : boolean;
  signal type_cast_1399_inst_req_1 : boolean;
  signal type_cast_1399_inst_ack_1 : boolean;
  signal type_cast_1395_inst_req_0 : boolean;
  signal if_stmt_1381_branch_ack_0 : boolean;
  signal if_stmt_1381_branch_ack_1 : boolean;
  signal phi_stmt_1230_req_1 : boolean;
  signal call_stmt_1306_call_ack_1 : boolean;
  signal call_stmt_1306_call_req_1 : boolean;
  signal do_while_stmt_1218_branch_ack_1 : boolean;
  signal type_cast_1395_inst_ack_1 : boolean;
  signal type_cast_1395_inst_req_1 : boolean;
  signal type_cast_1251_inst_req_0 : boolean;
  signal type_cast_1228_inst_ack_0 : boolean;
  signal type_cast_1346_inst_ack_0 : boolean;
  signal if_stmt_1381_branch_req_0 : boolean;
  signal type_cast_1228_inst_req_0 : boolean;
  signal type_cast_1346_inst_req_0 : boolean;
  signal phi_stmt_1230_req_0 : boolean;
  signal call_stmt_1306_call_ack_0 : boolean;
  signal W_row18x_x1x_xi_1329_delayed_2_0_1348_inst_ack_0 : boolean;
  signal call_stmt_1306_call_req_0 : boolean;
  signal W_row18x_x1x_xi_1329_delayed_2_0_1348_inst_req_0 : boolean;
  signal type_cast_1238_inst_ack_1 : boolean;
  signal type_cast_1238_inst_req_1 : boolean;
  signal do_while_stmt_1218_branch_ack_0 : boolean;
  signal type_cast_1346_inst_ack_1 : boolean;
  signal call_stmt_1192_call_req_0 : boolean;
  signal call_stmt_1192_call_ack_0 : boolean;
  signal call_stmt_1192_call_req_1 : boolean;
  signal call_stmt_1192_call_ack_1 : boolean;
  signal call_stmt_1194_call_req_0 : boolean;
  signal call_stmt_1194_call_ack_0 : boolean;
  signal call_stmt_1194_call_req_1 : boolean;
  signal call_stmt_1194_call_ack_1 : boolean;
  signal do_while_stmt_1218_branch_req_0 : boolean;
  signal phi_stmt_1220_req_0 : boolean;
  signal phi_stmt_1220_req_1 : boolean;
  signal phi_stmt_1220_ack_0 : boolean;
  signal W_iNsTr_2_1278_delayed_1_0_1293_inst_ack_0 : boolean;
  signal type_cast_1223_inst_req_0 : boolean;
  signal type_cast_1223_inst_ack_0 : boolean;
  signal type_cast_1223_inst_req_1 : boolean;
  signal type_cast_1223_inst_ack_1 : boolean;
  signal phi_stmt_1225_req_0 : boolean;
  signal phi_stmt_1225_req_1 : boolean;
  signal phi_stmt_1225_ack_0 : boolean;
  signal WPIPE_system_output_pipe_1401_inst_req_0 : boolean;
  signal WPIPE_system_output_pipe_1401_inst_ack_0 : boolean;
  signal WPIPE_system_output_pipe_1401_inst_req_1 : boolean;
  signal WPIPE_system_output_pipe_1401_inst_ack_1 : boolean;
  signal call_stmt_1405_call_req_0 : boolean;
  signal call_stmt_1405_call_ack_0 : boolean;
  signal call_stmt_1405_call_req_1 : boolean;
  signal call_stmt_1405_call_ack_1 : boolean;
  signal type_cast_1409_inst_req_0 : boolean;
  signal type_cast_1409_inst_ack_0 : boolean;
  signal type_cast_1409_inst_req_1 : boolean;
  signal type_cast_1409_inst_ack_1 : boolean;
  signal type_cast_1418_inst_req_0 : boolean;
  signal type_cast_1418_inst_ack_0 : boolean;
  signal type_cast_1418_inst_req_1 : boolean;
  signal type_cast_1418_inst_ack_1 : boolean;
  signal type_cast_1428_inst_req_0 : boolean;
  signal type_cast_1428_inst_ack_0 : boolean;
  signal type_cast_1428_inst_req_1 : boolean;
  signal type_cast_1428_inst_ack_1 : boolean;
  signal type_cast_1438_inst_req_0 : boolean;
  signal type_cast_1438_inst_ack_0 : boolean;
  signal type_cast_1438_inst_req_1 : boolean;
  signal type_cast_1438_inst_ack_1 : boolean;
  signal type_cast_1448_inst_req_0 : boolean;
  signal type_cast_1448_inst_ack_0 : boolean;
  signal type_cast_1448_inst_req_1 : boolean;
  signal type_cast_1448_inst_ack_1 : boolean;
  signal type_cast_1458_inst_req_0 : boolean;
  signal type_cast_1458_inst_ack_0 : boolean;
  signal type_cast_1458_inst_req_1 : boolean;
  signal type_cast_1458_inst_ack_1 : boolean;
  signal type_cast_1468_inst_req_0 : boolean;
  signal type_cast_1468_inst_ack_0 : boolean;
  signal type_cast_1468_inst_req_1 : boolean;
  signal type_cast_1468_inst_ack_1 : boolean;
  signal type_cast_1478_inst_req_0 : boolean;
  signal type_cast_1478_inst_ack_0 : boolean;
  signal type_cast_1478_inst_req_1 : boolean;
  signal type_cast_1478_inst_ack_1 : boolean;
  signal type_cast_1488_inst_req_0 : boolean;
  signal type_cast_1488_inst_ack_0 : boolean;
  signal type_cast_1488_inst_req_1 : boolean;
  signal type_cast_1488_inst_ack_1 : boolean;
  signal WPIPE_system_output_pipe_1490_inst_req_0 : boolean;
  signal WPIPE_system_output_pipe_1490_inst_ack_0 : boolean;
  signal WPIPE_system_output_pipe_1490_inst_req_1 : boolean;
  signal WPIPE_system_output_pipe_1490_inst_ack_1 : boolean;
  signal WPIPE_system_output_pipe_1493_inst_req_0 : boolean;
  signal WPIPE_system_output_pipe_1493_inst_ack_0 : boolean;
  signal WPIPE_system_output_pipe_1493_inst_req_1 : boolean;
  signal WPIPE_system_output_pipe_1493_inst_ack_1 : boolean;
  signal WPIPE_system_output_pipe_1496_inst_req_0 : boolean;
  signal WPIPE_system_output_pipe_1496_inst_ack_0 : boolean;
  signal WPIPE_system_output_pipe_1496_inst_req_1 : boolean;
  signal WPIPE_system_output_pipe_1496_inst_ack_1 : boolean;
  signal WPIPE_system_output_pipe_1499_inst_req_0 : boolean;
  signal WPIPE_system_output_pipe_1499_inst_ack_0 : boolean;
  signal WPIPE_system_output_pipe_1499_inst_req_1 : boolean;
  signal WPIPE_system_output_pipe_1499_inst_ack_1 : boolean;
  signal WPIPE_system_output_pipe_1502_inst_req_0 : boolean;
  signal WPIPE_system_output_pipe_1502_inst_ack_0 : boolean;
  signal WPIPE_system_output_pipe_1502_inst_req_1 : boolean;
  signal WPIPE_system_output_pipe_1502_inst_ack_1 : boolean;
  signal WPIPE_system_output_pipe_1505_inst_req_0 : boolean;
  signal WPIPE_system_output_pipe_1505_inst_ack_0 : boolean;
  signal WPIPE_system_output_pipe_1505_inst_req_1 : boolean;
  signal WPIPE_system_output_pipe_1505_inst_ack_1 : boolean;
  signal WPIPE_system_output_pipe_1508_inst_req_0 : boolean;
  signal WPIPE_system_output_pipe_1508_inst_ack_0 : boolean;
  signal WPIPE_system_output_pipe_1508_inst_req_1 : boolean;
  signal WPIPE_system_output_pipe_1508_inst_ack_1 : boolean;
  signal WPIPE_system_output_pipe_1511_inst_req_0 : boolean;
  signal WPIPE_system_output_pipe_1511_inst_ack_0 : boolean;
  signal WPIPE_system_output_pipe_1511_inst_req_1 : boolean;
  signal WPIPE_system_output_pipe_1511_inst_ack_1 : boolean;
  signal call_stmt_1514_call_req_0 : boolean;
  signal call_stmt_1514_call_ack_0 : boolean;
  signal call_stmt_1514_call_req_1 : boolean;
  signal call_stmt_1514_call_ack_1 : boolean;
  signal type_cast_1389_inst_req_0 : boolean;
  signal type_cast_1389_inst_ack_0 : boolean;
  signal type_cast_1389_inst_req_1 : boolean;
  signal type_cast_1389_inst_ack_1 : boolean;
  signal phi_stmt_1386_req_0 : boolean;
  signal phi_stmt_1386_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "systemTOP_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  systemTOP_CP_2045_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "systemTOP_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= systemTOP_CP_2045_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= systemTOP_CP_2045_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= systemTOP_CP_2045_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  systemTOP_CP_2045: Block -- control-path 
    signal systemTOP_CP_2045_elements: BooleanArray(208 downto 0);
    -- 
  begin -- 
    systemTOP_CP_2045_elements(0) <= systemTOP_CP_2045_start;
    systemTOP_CP_2045_symbol <= systemTOP_CP_2045_elements(204);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0:  members (17) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1191/$entry
      -- CP-element group 0: 	 branch_block_stmt_1191/branch_block_stmt_1191__entry__
      -- CP-element group 0: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194__entry__
      -- CP-element group 0: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/$entry
      -- CP-element group 0: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1192_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1192_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1192_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1192_Sample/crr
      -- CP-element group 0: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1192_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1192_Update/ccr
      -- CP-element group 0: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1194_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1194_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1194_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1194_Sample/crr
      -- CP-element group 0: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1194_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1194_Update/ccr
      -- 
    crr_2077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(0), ack => call_stmt_1192_call_req_0); -- 
    ccr_2082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(0), ack => call_stmt_1192_call_req_1); -- 
    crr_2091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(0), ack => call_stmt_1194_call_req_0); -- 
    ccr_2096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(0), ack => call_stmt_1194_call_req_1); -- 
    -- CP-element group 1:  branch  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	142 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	143 
    -- CP-element group 1: 	144 
    -- CP-element group 1:  members (9) 
      -- CP-element group 1: 	 branch_block_stmt_1191/if_stmt_1381_dead_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1191/if_stmt_1381_eval_test/$exit
      -- CP-element group 1: 	 branch_block_stmt_1191/if_stmt_1381_else_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1191/if_stmt_1381_if_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1191/if_stmt_1381_eval_test/$entry
      -- CP-element group 1: 	 branch_block_stmt_1191/R_whilex_xbodyx_xi_maxPool3Dx_xexit_taken_1382_place
      -- CP-element group 1: 	 branch_block_stmt_1191/if_stmt_1381_eval_test/branch_req
      -- CP-element group 1: 	 branch_block_stmt_1191/do_while_stmt_1218__exit__
      -- CP-element group 1: 	 branch_block_stmt_1191/if_stmt_1381__entry__
      -- 
    branch_req_2437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(1), ack => if_stmt_1381_branch_req_0); -- 
    systemTOP_CP_2045_elements(1) <= systemTOP_CP_2045_elements(142);
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1192_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1192_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1192_Sample/cra
      -- 
    cra_2078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1192_call_ack_0, ack => systemTOP_CP_2045_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1192_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1192_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1192_Update/cca
      -- 
    cca_2083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1192_call_ack_1, ack => systemTOP_CP_2045_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1194_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1194_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1194_Sample/cra
      -- 
    cra_2092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1194_call_ack_0, ack => systemTOP_CP_2045_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1194_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1194_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/call_stmt_1194_Update/cca
      -- 
    cca_2097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1194_call_ack_1, ack => systemTOP_CP_2045_elements(5)); -- 
    -- CP-element group 6:  join  transition  place  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: 	3 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (10) 
      -- CP-element group 6: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194__exit__
      -- CP-element group 6: 	 branch_block_stmt_1191/entry_whilex_xbodyx_xi
      -- CP-element group 6: 	 branch_block_stmt_1191/merge_stmt_1196__exit__
      -- CP-element group 6: 	 branch_block_stmt_1191/do_while_stmt_1218__entry__
      -- CP-element group 6: 	 branch_block_stmt_1191/call_stmt_1192_to_call_stmt_1194/$exit
      -- CP-element group 6: 	 branch_block_stmt_1191/entry_whilex_xbodyx_xi_PhiReq/$entry
      -- CP-element group 6: 	 branch_block_stmt_1191/entry_whilex_xbodyx_xi_PhiReq/$exit
      -- CP-element group 6: 	 branch_block_stmt_1191/merge_stmt_1196_PhiReqMerge
      -- CP-element group 6: 	 branch_block_stmt_1191/merge_stmt_1196_PhiAck/$entry
      -- CP-element group 6: 	 branch_block_stmt_1191/merge_stmt_1196_PhiAck/$exit
      -- 
    systemTOP_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "systemTOP_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(5) & systemTOP_CP_2045_elements(3);
      gj_systemTOP_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_1191/do_while_stmt_1218/$entry
      -- CP-element group 7: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218__entry__
      -- 
    systemTOP_CP_2045_elements(7) <= systemTOP_CP_2045_elements(6);
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	142 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218__exit__
      -- 
    -- Element group systemTOP_CP_2045_elements(8) is bound as output of CP function.
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1191/do_while_stmt_1218/loop_back
      -- 
    -- Element group systemTOP_CP_2045_elements(9) is bound as output of CP function.
    -- CP-element group 10:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	140 
    -- CP-element group 10: 	141 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1191/do_while_stmt_1218/loop_taken/$entry
      -- CP-element group 10: 	 branch_block_stmt_1191/do_while_stmt_1218/loop_exit/$entry
      -- CP-element group 10: 	 branch_block_stmt_1191/do_while_stmt_1218/condition_done
      -- 
    systemTOP_CP_2045_elements(10) <= systemTOP_CP_2045_elements(15);
    -- CP-element group 11:  branch  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	139 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1191/do_while_stmt_1218/loop_body_done
      -- 
    systemTOP_CP_2045_elements(11) <= systemTOP_CP_2045_elements(139);
    -- CP-element group 12:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	45 
    -- CP-element group 12: 	87 
    -- CP-element group 12: 	66 
    -- CP-element group 12: 	26 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/back_edge_to_loop_body
      -- 
    systemTOP_CP_2045_elements(12) <= systemTOP_CP_2045_elements(9);
    -- CP-element group 13:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	47 
    -- CP-element group 13: 	89 
    -- CP-element group 13: 	68 
    -- CP-element group 13: 	28 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/first_time_through_loop_body
      -- 
    systemTOP_CP_2045_elements(13) <= systemTOP_CP_2045_elements(7);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	42 
    -- CP-element group 14: 	138 
    -- CP-element group 14: 	60 
    -- CP-element group 14: 	82 
    -- CP-element group 14: 	81 
    -- CP-element group 14: 	61 
    -- CP-element group 14: 	41 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	21 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/$entry
      -- CP-element group 14: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/loop_body_start
      -- 
    -- Element group systemTOP_CP_2045_elements(14) is bound as output of CP function.
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	133 
    -- CP-element group 15: 	137 
    -- CP-element group 15: 	138 
    -- CP-element group 15: 	19 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/condition_evaluated
      -- 
    condition_evaluated_2112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(15), ack => do_while_stmt_1218_branch_req_0); -- 
    systemTOP_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "systemTOP_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(133) & systemTOP_CP_2045_elements(137) & systemTOP_CP_2045_elements(138) & systemTOP_CP_2045_elements(19);
      gj_systemTOP_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	60 
    -- CP-element group 16: 	81 
    -- CP-element group 16: 	41 
    -- CP-element group 16: 	20 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	19 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	83 
    -- CP-element group 16: 	62 
    -- CP-element group 16: 	22 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/aggregated_phi_sample_req
      -- CP-element group 16: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1225_sample_start__ps
      -- 
    systemTOP_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "systemTOP_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(60) & systemTOP_CP_2045_elements(81) & systemTOP_CP_2045_elements(41) & systemTOP_CP_2045_elements(20) & systemTOP_CP_2045_elements(19);
      gj_systemTOP_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	43 
    -- CP-element group 17: 	84 
    -- CP-element group 17: 	63 
    -- CP-element group 17: 	23 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	123 
    -- CP-element group 17: 	127 
    -- CP-element group 17: 	131 
    -- CP-element group 17: 	135 
    -- CP-element group 17: 	139 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	60 
    -- CP-element group 17: 	81 
    -- CP-element group 17: 	41 
    -- CP-element group 17: 	20 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1235_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1230_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/aggregated_phi_sample_ack
      -- CP-element group 17: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1220_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1225_sample_completed_
      -- 
    systemTOP_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "systemTOP_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(43) & systemTOP_CP_2045_elements(84) & systemTOP_CP_2045_elements(63) & systemTOP_CP_2045_elements(23);
      gj_systemTOP_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	42 
    -- CP-element group 18: 	82 
    -- CP-element group 18: 	61 
    -- CP-element group 18: 	21 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	85 
    -- CP-element group 18: 	64 
    -- CP-element group 18: 	24 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/aggregated_phi_update_req
      -- CP-element group 18: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1225_update_start__ps
      -- 
    systemTOP_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "systemTOP_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(42) & systemTOP_CP_2045_elements(82) & systemTOP_CP_2045_elements(61) & systemTOP_CP_2045_elements(21);
      gj_systemTOP_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	44 
    -- CP-element group 19: 	86 
    -- CP-element group 19: 	65 
    -- CP-element group 19: 	25 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	16 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/aggregated_phi_update_ack
      -- 
    systemTOP_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "systemTOP_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(44) & systemTOP_CP_2045_elements(86) & systemTOP_CP_2045_elements(65) & systemTOP_CP_2045_elements(25);
      gj_systemTOP_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	17 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1220_sample_start_
      -- 
    systemTOP_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "systemTOP_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(14) & systemTOP_CP_2045_elements(17);
      gj_systemTOP_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	14 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	116 
    -- CP-element group 21: 	25 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	18 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1220_update_start_
      -- 
    systemTOP_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "systemTOP_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(14) & systemTOP_CP_2045_elements(116) & systemTOP_CP_2045_elements(25);
      gj_systemTOP_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	16 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1220_sample_start__ps
      -- 
    systemTOP_CP_2045_elements(22) <= systemTOP_CP_2045_elements(16);
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	17 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1220_sample_completed__ps
      -- 
    -- Element group systemTOP_CP_2045_elements(23) is bound as output of CP function.
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	18 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1220_update_start__ps
      -- 
    systemTOP_CP_2045_elements(24) <= systemTOP_CP_2045_elements(18);
    -- CP-element group 25:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	114 
    -- CP-element group 25: 	19 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	21 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1220_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1220_update_completed__ps
      -- 
    -- Element group systemTOP_CP_2045_elements(25) is bound as output of CP function.
    -- CP-element group 26:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	12 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1220_loopback_trigger
      -- 
    systemTOP_CP_2045_elements(26) <= systemTOP_CP_2045_elements(12);
    -- CP-element group 27:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1220_loopback_sample_req
      -- CP-element group 27: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1220_loopback_sample_req_ps
      -- 
    phi_stmt_1220_loopback_sample_req_2127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1220_loopback_sample_req_2127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(27), ack => phi_stmt_1220_req_0); -- 
    -- Element group systemTOP_CP_2045_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	13 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1220_entry_trigger
      -- 
    systemTOP_CP_2045_elements(28) <= systemTOP_CP_2045_elements(13);
    -- CP-element group 29:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1220_entry_sample_req
      -- CP-element group 29: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1220_entry_sample_req_ps
      -- 
    phi_stmt_1220_entry_sample_req_2130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1220_entry_sample_req_2130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(29), ack => phi_stmt_1220_req_1); -- 
    -- Element group systemTOP_CP_2045_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1220_phi_mux_ack
      -- CP-element group 30: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1220_phi_mux_ack_ps
      -- 
    phi_stmt_1220_phi_mux_ack_2133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1220_ack_0, ack => systemTOP_CP_2045_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1223_sample_start__ps
      -- 
    -- Element group systemTOP_CP_2045_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1223_update_start__ps
      -- 
    -- Element group systemTOP_CP_2045_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	35 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1223_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1223_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1223_Sample/rr
      -- 
    rr_2146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(33), ack => type_cast_1223_inst_req_0); -- 
    systemTOP_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "systemTOP_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(31) & systemTOP_CP_2045_elements(35);
      gj_systemTOP_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1223_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1223_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1223_Update/cr
      -- 
    cr_2151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(34), ack => type_cast_1223_inst_req_1); -- 
    systemTOP_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "systemTOP_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(32) & systemTOP_CP_2045_elements(36);
      gj_systemTOP_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	33 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1223_sample_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1223_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1223_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1223_Sample/ra
      -- 
    ra_2147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1223_inst_ack_0, ack => systemTOP_CP_2045_elements(35)); -- 
    -- CP-element group 36:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	34 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1223_update_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1223_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1223_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1223_Update/ca
      -- 
    ca_2152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1223_inst_ack_1, ack => systemTOP_CP_2045_elements(36)); -- 
    -- CP-element group 37:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_iNsTr_2_at_entry_1224_sample_start__ps
      -- CP-element group 37: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_iNsTr_2_at_entry_1224_sample_completed__ps
      -- CP-element group 37: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_iNsTr_2_at_entry_1224_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_iNsTr_2_at_entry_1224_sample_completed_
      -- 
    -- Element group systemTOP_CP_2045_elements(37) is bound as output of CP function.
    -- CP-element group 38:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_iNsTr_2_at_entry_1224_update_start__ps
      -- CP-element group 38: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_iNsTr_2_at_entry_1224_update_start_
      -- 
    -- Element group systemTOP_CP_2045_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	40 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_iNsTr_2_at_entry_1224_update_completed__ps
      -- 
    systemTOP_CP_2045_elements(39) <= systemTOP_CP_2045_elements(40);
    -- CP-element group 40:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	39 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_iNsTr_2_at_entry_1224_update_completed_
      -- 
    -- Element group systemTOP_CP_2045_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => systemTOP_CP_2045_elements(38), ack => systemTOP_CP_2045_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	14 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	133 
    -- CP-element group 41: 	137 
    -- CP-element group 41: 	17 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	16 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1225_sample_start_
      -- 
    systemTOP_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "systemTOP_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(14) & systemTOP_CP_2045_elements(133) & systemTOP_CP_2045_elements(137) & systemTOP_CP_2045_elements(17);
      gj_systemTOP_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  join  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	14 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	112 
    -- CP-element group 42: 	44 
    -- CP-element group 42: 	136 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	18 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1225_update_start_
      -- 
    systemTOP_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "systemTOP_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(14) & systemTOP_CP_2045_elements(112) & systemTOP_CP_2045_elements(44) & systemTOP_CP_2045_elements(136);
      gj_systemTOP_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  join  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	17 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1225_sample_completed__ps
      -- 
    -- Element group systemTOP_CP_2045_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	110 
    -- CP-element group 44: 	134 
    -- CP-element group 44: 	19 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1225_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1225_update_completed__ps
      -- 
    -- Element group systemTOP_CP_2045_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	12 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1225_loopback_trigger
      -- 
    systemTOP_CP_2045_elements(45) <= systemTOP_CP_2045_elements(12);
    -- CP-element group 46:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1225_loopback_sample_req
      -- CP-element group 46: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1225_loopback_sample_req_ps
      -- 
    phi_stmt_1225_loopback_sample_req_2171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1225_loopback_sample_req_2171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(46), ack => phi_stmt_1225_req_0); -- 
    -- Element group systemTOP_CP_2045_elements(46) is bound as output of CP function.
    -- CP-element group 47:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	13 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1225_entry_trigger
      -- 
    systemTOP_CP_2045_elements(47) <= systemTOP_CP_2045_elements(13);
    -- CP-element group 48:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1225_entry_sample_req
      -- CP-element group 48: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1225_entry_sample_req_ps
      -- 
    phi_stmt_1225_entry_sample_req_2174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1225_entry_sample_req_2174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(48), ack => phi_stmt_1225_req_1); -- 
    -- Element group systemTOP_CP_2045_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1225_phi_mux_ack
      -- CP-element group 49: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1225_phi_mux_ack_ps
      -- 
    phi_stmt_1225_phi_mux_ack_2177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1225_ack_0, ack => systemTOP_CP_2045_elements(49)); -- 
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1228_sample_start__ps
      -- 
    -- Element group systemTOP_CP_2045_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1228_update_start__ps
      -- 
    -- Element group systemTOP_CP_2045_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1228_Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1228_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1228_sample_start_
      -- 
    rr_2190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(52), ack => type_cast_1228_inst_req_0); -- 
    systemTOP_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "systemTOP_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(50) & systemTOP_CP_2045_elements(54);
      gj_systemTOP_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	55 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1228_Update/cr
      -- CP-element group 53: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1228_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1228_update_start_
      -- 
    cr_2195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(53), ack => type_cast_1228_inst_req_1); -- 
    systemTOP_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "systemTOP_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(51) & systemTOP_CP_2045_elements(55);
      gj_systemTOP_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	52 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1228_Sample/ra
      -- CP-element group 54: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1228_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1228_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1228_sample_completed__ps
      -- 
    ra_2191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1228_inst_ack_0, ack => systemTOP_CP_2045_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: marked-successors 
    -- CP-element group 55: 	53 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1228_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1228_Update/ca
      -- CP-element group 55: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1228_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1228_update_completed__ps
      -- 
    ca_2196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1228_inst_ack_1, ack => systemTOP_CP_2045_elements(55)); -- 
    -- CP-element group 56:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_row18x_x1x_xi_at_entry_1229_sample_completed__ps
      -- CP-element group 56: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_row18x_x1x_xi_at_entry_1229_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_row18x_x1x_xi_at_entry_1229_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_row18x_x1x_xi_at_entry_1229_sample_start__ps
      -- 
    -- Element group systemTOP_CP_2045_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_row18x_x1x_xi_at_entry_1229_update_start__ps
      -- CP-element group 57: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_row18x_x1x_xi_at_entry_1229_update_start_
      -- 
    -- Element group systemTOP_CP_2045_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_row18x_x1x_xi_at_entry_1229_update_completed__ps
      -- 
    systemTOP_CP_2045_elements(58) <= systemTOP_CP_2045_elements(59);
    -- CP-element group 59:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	58 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_row18x_x1x_xi_at_entry_1229_update_completed_
      -- 
    -- Element group systemTOP_CP_2045_elements(59) is a control-delay.
    cp_element_59_delay: control_delay_element  generic map(name => " 59_delay", delay_value => 1)  port map(req => systemTOP_CP_2045_elements(57), ack => systemTOP_CP_2045_elements(59), clk => clk, reset =>reset);
    -- CP-element group 60:  join  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	14 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	125 
    -- CP-element group 60: 	129 
    -- CP-element group 60: 	17 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	16 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1230_sample_start_
      -- 
    systemTOP_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "systemTOP_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(14) & systemTOP_CP_2045_elements(125) & systemTOP_CP_2045_elements(129) & systemTOP_CP_2045_elements(17);
      gj_systemTOP_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  join  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	14 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	108 
    -- CP-element group 61: 	128 
    -- CP-element group 61: 	65 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	18 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1230_update_start_
      -- 
    systemTOP_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "systemTOP_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(14) & systemTOP_CP_2045_elements(108) & systemTOP_CP_2045_elements(128) & systemTOP_CP_2045_elements(65);
      gj_systemTOP_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	16 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1230_sample_start__ps
      -- 
    systemTOP_CP_2045_elements(62) <= systemTOP_CP_2045_elements(16);
    -- CP-element group 63:  join  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	17 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1230_sample_completed__ps
      -- 
    -- Element group systemTOP_CP_2045_elements(63) is bound as output of CP function.
    -- CP-element group 64:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	18 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1230_update_start__ps
      -- 
    systemTOP_CP_2045_elements(64) <= systemTOP_CP_2045_elements(18);
    -- CP-element group 65:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	106 
    -- CP-element group 65: 	126 
    -- CP-element group 65: 	19 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	61 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1230_update_completed__ps
      -- CP-element group 65: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1230_update_completed_
      -- 
    -- Element group systemTOP_CP_2045_elements(65) is bound as output of CP function.
    -- CP-element group 66:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	12 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1230_loopback_trigger
      -- 
    systemTOP_CP_2045_elements(66) <= systemTOP_CP_2045_elements(12);
    -- CP-element group 67:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1230_loopback_sample_req_ps
      -- CP-element group 67: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1230_loopback_sample_req
      -- 
    phi_stmt_1230_loopback_sample_req_2215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1230_loopback_sample_req_2215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(67), ack => phi_stmt_1230_req_0); -- 
    -- Element group systemTOP_CP_2045_elements(67) is bound as output of CP function.
    -- CP-element group 68:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	13 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1230_entry_trigger
      -- 
    systemTOP_CP_2045_elements(68) <= systemTOP_CP_2045_elements(13);
    -- CP-element group 69:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1230_entry_sample_req_ps
      -- CP-element group 69: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1230_entry_sample_req
      -- 
    phi_stmt_1230_entry_sample_req_2218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1230_entry_sample_req_2218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(69), ack => phi_stmt_1230_req_1); -- 
    -- Element group systemTOP_CP_2045_elements(69) is bound as output of CP function.
    -- CP-element group 70:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1230_phi_mux_ack_ps
      -- CP-element group 70: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1230_phi_mux_ack
      -- 
    phi_stmt_1230_phi_mux_ack_2221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1230_ack_0, ack => systemTOP_CP_2045_elements(70)); -- 
    -- CP-element group 71:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1233_sample_start__ps
      -- 
    -- Element group systemTOP_CP_2045_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1233_update_start__ps
      -- 
    -- Element group systemTOP_CP_2045_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	75 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1233_Sample/rr
      -- CP-element group 73: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1233_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1233_sample_start_
      -- 
    rr_2234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(73), ack => type_cast_1233_inst_req_0); -- 
    systemTOP_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "systemTOP_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(71) & systemTOP_CP_2045_elements(75);
      gj_systemTOP_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1233_Update/cr
      -- CP-element group 74: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1233_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1233_update_start_
      -- 
    cr_2239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(74), ack => type_cast_1233_inst_req_1); -- 
    systemTOP_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "systemTOP_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(72) & systemTOP_CP_2045_elements(76);
      gj_systemTOP_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	73 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1233_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1233_sample_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1233_Sample/ra
      -- CP-element group 75: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1233_sample_completed_
      -- 
    ra_2235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1233_inst_ack_0, ack => systemTOP_CP_2045_elements(75)); -- 
    -- CP-element group 76:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	74 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1233_Update/ca
      -- CP-element group 76: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1233_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1233_update_completed__ps
      -- CP-element group 76: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1233_update_completed_
      -- 
    ca_2240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1233_inst_ack_1, ack => systemTOP_CP_2045_elements(76)); -- 
    -- CP-element group 77:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (4) 
      -- CP-element group 77: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_colx_x1x_xi_at_entry_1234_sample_start__ps
      -- CP-element group 77: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_colx_x1x_xi_at_entry_1234_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_colx_x1x_xi_at_entry_1234_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_colx_x1x_xi_at_entry_1234_sample_completed__ps
      -- 
    -- Element group systemTOP_CP_2045_elements(77) is bound as output of CP function.
    -- CP-element group 78:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_colx_x1x_xi_at_entry_1234_update_start_
      -- CP-element group 78: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_colx_x1x_xi_at_entry_1234_update_start__ps
      -- 
    -- Element group systemTOP_CP_2045_elements(78) is bound as output of CP function.
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_colx_x1x_xi_at_entry_1234_update_completed__ps
      -- 
    systemTOP_CP_2045_elements(79) <= systemTOP_CP_2045_elements(80);
    -- CP-element group 80:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	79 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_colx_x1x_xi_at_entry_1234_update_completed_
      -- 
    -- Element group systemTOP_CP_2045_elements(80) is a control-delay.
    cp_element_80_delay: control_delay_element  generic map(name => " 80_delay", delay_value => 1)  port map(req => systemTOP_CP_2045_elements(78), ack => systemTOP_CP_2045_elements(80), clk => clk, reset =>reset);
    -- CP-element group 81:  join  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	14 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	17 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	16 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1235_sample_start_
      -- 
    systemTOP_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "systemTOP_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(14) & systemTOP_CP_2045_elements(17);
      gj_systemTOP_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  join  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	14 
    -- CP-element group 82: marked-predecessors 
    -- CP-element group 82: 	104 
    -- CP-element group 82: 	124 
    -- CP-element group 82: 	86 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	18 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1235_update_start_
      -- 
    systemTOP_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "systemTOP_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(14) & systemTOP_CP_2045_elements(104) & systemTOP_CP_2045_elements(124) & systemTOP_CP_2045_elements(86);
      gj_systemTOP_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	16 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1235_sample_start__ps
      -- 
    systemTOP_CP_2045_elements(83) <= systemTOP_CP_2045_elements(16);
    -- CP-element group 84:  join  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	17 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1235_sample_completed__ps
      -- 
    -- Element group systemTOP_CP_2045_elements(84) is bound as output of CP function.
    -- CP-element group 85:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	18 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1235_update_start__ps
      -- 
    systemTOP_CP_2045_elements(85) <= systemTOP_CP_2045_elements(18);
    -- CP-element group 86:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	102 
    -- CP-element group 86: 	122 
    -- CP-element group 86: 	19 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	82 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1235_update_completed__ps
      -- CP-element group 86: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1235_update_completed_
      -- 
    -- Element group systemTOP_CP_2045_elements(86) is bound as output of CP function.
    -- CP-element group 87:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	12 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1235_loopback_trigger
      -- 
    systemTOP_CP_2045_elements(87) <= systemTOP_CP_2045_elements(12);
    -- CP-element group 88:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1235_loopback_sample_req
      -- CP-element group 88: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1235_loopback_sample_req_ps
      -- 
    phi_stmt_1235_loopback_sample_req_2259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1235_loopback_sample_req_2259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(88), ack => phi_stmt_1235_req_0); -- 
    -- Element group systemTOP_CP_2045_elements(88) is bound as output of CP function.
    -- CP-element group 89:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	13 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1235_entry_trigger
      -- 
    systemTOP_CP_2045_elements(89) <= systemTOP_CP_2045_elements(13);
    -- CP-element group 90:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1235_entry_sample_req
      -- CP-element group 90: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1235_entry_sample_req_ps
      -- 
    phi_stmt_1235_entry_sample_req_2262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1235_entry_sample_req_2262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(90), ack => phi_stmt_1235_req_1); -- 
    -- Element group systemTOP_CP_2045_elements(90) is bound as output of CP function.
    -- CP-element group 91:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1235_phi_mux_ack
      -- CP-element group 91: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/phi_stmt_1235_phi_mux_ack_ps
      -- 
    phi_stmt_1235_phi_mux_ack_2265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1235_ack_0, ack => systemTOP_CP_2045_elements(91)); -- 
    -- CP-element group 92:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1238_sample_start__ps
      -- 
    -- Element group systemTOP_CP_2045_elements(92) is bound as output of CP function.
    -- CP-element group 93:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1238_update_start__ps
      -- 
    -- Element group systemTOP_CP_2045_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	96 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1238_Sample/rr
      -- CP-element group 94: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1238_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1238_Sample/$entry
      -- 
    rr_2278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(94), ack => type_cast_1238_inst_req_0); -- 
    systemTOP_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "systemTOP_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(92) & systemTOP_CP_2045_elements(96);
      gj_systemTOP_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	97 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1238_update_start_
      -- CP-element group 95: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1238_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1238_Update/cr
      -- 
    cr_2283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(95), ack => type_cast_1238_inst_req_1); -- 
    systemTOP_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "systemTOP_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(93) & systemTOP_CP_2045_elements(97);
      gj_systemTOP_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	94 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1238_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1238_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1238_sample_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1238_Sample/ra
      -- 
    ra_2279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_0, ack => systemTOP_CP_2045_elements(96)); -- 
    -- CP-element group 97:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: marked-successors 
    -- CP-element group 97: 	95 
    -- CP-element group 97:  members (4) 
      -- CP-element group 97: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1238_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1238_update_completed__ps
      -- CP-element group 97: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1238_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1238_Update/$exit
      -- 
    ca_2284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_1, ack => systemTOP_CP_2045_elements(97)); -- 
    -- CP-element group 98:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (4) 
      -- CP-element group 98: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_chlx_x0x_xi_at_entry_1239_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_chlx_x0x_xi_at_entry_1239_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_chlx_x0x_xi_at_entry_1239_sample_completed__ps
      -- CP-element group 98: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_chlx_x0x_xi_at_entry_1239_sample_start__ps
      -- 
    -- Element group systemTOP_CP_2045_elements(98) is bound as output of CP function.
    -- CP-element group 99:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_chlx_x0x_xi_at_entry_1239_update_start_
      -- CP-element group 99: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_chlx_x0x_xi_at_entry_1239_update_start__ps
      -- 
    -- Element group systemTOP_CP_2045_elements(99) is bound as output of CP function.
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	101 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_chlx_x0x_xi_at_entry_1239_update_completed__ps
      -- 
    systemTOP_CP_2045_elements(100) <= systemTOP_CP_2045_elements(101);
    -- CP-element group 101:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	100 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/R_chlx_x0x_xi_at_entry_1239_update_completed_
      -- 
    -- Element group systemTOP_CP_2045_elements(101) is a control-delay.
    cp_element_101_delay: control_delay_element  generic map(name => " 101_delay", delay_value => 1)  port map(req => systemTOP_CP_2045_elements(99), ack => systemTOP_CP_2045_elements(101), clk => clk, reset =>reset);
    -- CP-element group 102:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	86 
    -- CP-element group 102: marked-predecessors 
    -- CP-element group 102: 	104 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1243_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1243_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1243_sample_start_
      -- 
    rr_2301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(102), ack => type_cast_1243_inst_req_0); -- 
    systemTOP_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(86) & systemTOP_CP_2045_elements(104);
      gj_systemTOP_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: marked-predecessors 
    -- CP-element group 103: 	105 
    -- CP-element group 103: 	120 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1243_Update/cr
      -- CP-element group 103: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1243_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1243_update_start_
      -- 
    cr_2306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(103), ack => type_cast_1243_inst_req_1); -- 
    systemTOP_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(105) & systemTOP_CP_2045_elements(120);
      gj_systemTOP_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104: marked-successors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	82 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1243_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1243_Sample/ra
      -- CP-element group 104: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1243_Sample/$exit
      -- 
    ra_2302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1243_inst_ack_0, ack => systemTOP_CP_2045_elements(104)); -- 
    -- CP-element group 105:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	118 
    -- CP-element group 105: marked-successors 
    -- CP-element group 105: 	103 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1243_Update/ca
      -- CP-element group 105: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1243_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1243_Update/$exit
      -- 
    ca_2307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1243_inst_ack_1, ack => systemTOP_CP_2045_elements(105)); -- 
    -- CP-element group 106:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	65 
    -- CP-element group 106: marked-predecessors 
    -- CP-element group 106: 	108 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1247_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1247_Sample/rr
      -- CP-element group 106: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1247_Sample/$entry
      -- 
    rr_2315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(106), ack => type_cast_1247_inst_req_0); -- 
    systemTOP_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(65) & systemTOP_CP_2045_elements(108);
      gj_systemTOP_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: marked-predecessors 
    -- CP-element group 107: 	109 
    -- CP-element group 107: 	120 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1247_Update/cr
      -- CP-element group 107: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1247_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1247_update_start_
      -- 
    cr_2320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(107), ack => type_cast_1247_inst_req_1); -- 
    systemTOP_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(109) & systemTOP_CP_2045_elements(120);
      gj_systemTOP_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108: marked-successors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	61 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1247_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1247_Sample/ra
      -- CP-element group 108: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1247_Sample/$exit
      -- 
    ra_2316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1247_inst_ack_0, ack => systemTOP_CP_2045_elements(108)); -- 
    -- CP-element group 109:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	118 
    -- CP-element group 109: marked-successors 
    -- CP-element group 109: 	107 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1247_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1247_Update/ca
      -- CP-element group 109: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1247_update_completed_
      -- 
    ca_2321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1247_inst_ack_1, ack => systemTOP_CP_2045_elements(109)); -- 
    -- CP-element group 110:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	44 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	112 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1251_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1251_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1251_Sample/rr
      -- 
    rr_2329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(110), ack => type_cast_1251_inst_req_0); -- 
    systemTOP_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(44) & systemTOP_CP_2045_elements(112);
      gj_systemTOP_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: marked-predecessors 
    -- CP-element group 111: 	113 
    -- CP-element group 111: 	120 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1251_update_start_
      -- CP-element group 111: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1251_Update/cr
      -- CP-element group 111: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1251_Update/$entry
      -- 
    cr_2334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(111), ack => type_cast_1251_inst_req_1); -- 
    systemTOP_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(113) & systemTOP_CP_2045_elements(120);
      gj_systemTOP_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: marked-successors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: 	42 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1251_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1251_Sample/ra
      -- CP-element group 112: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1251_Sample/$exit
      -- 
    ra_2330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1251_inst_ack_0, ack => systemTOP_CP_2045_elements(112)); -- 
    -- CP-element group 113:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	118 
    -- CP-element group 113: marked-successors 
    -- CP-element group 113: 	111 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1251_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1251_Update/ca
      -- CP-element group 113: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1251_Update/$exit
      -- 
    ca_2335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1251_inst_ack_1, ack => systemTOP_CP_2045_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	25 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	116 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1295_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1295_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1295_Sample/req
      -- 
    req_2343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(114), ack => W_iNsTr_2_1278_delayed_1_0_1293_inst_req_0); -- 
    systemTOP_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(25) & systemTOP_CP_2045_elements(116);
      gj_systemTOP_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: marked-predecessors 
    -- CP-element group 115: 	117 
    -- CP-element group 115: 	120 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1295_Update/req
      -- CP-element group 115: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1295_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1295_update_start_
      -- 
    req_2348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(115), ack => W_iNsTr_2_1278_delayed_1_0_1293_inst_req_1); -- 
    systemTOP_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(117) & systemTOP_CP_2045_elements(120);
      gj_systemTOP_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: marked-successors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: 	21 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1295_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1295_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1295_Sample/ack
      -- 
    ack_2344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iNsTr_2_1278_delayed_1_0_1293_inst_ack_0, ack => systemTOP_CP_2045_elements(116)); -- 
    -- CP-element group 117:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	115 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1295_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1295_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1295_Update/ack
      -- 
    ack_2349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iNsTr_2_1278_delayed_1_0_1293_inst_ack_1, ack => systemTOP_CP_2045_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	105 
    -- CP-element group 118: 	109 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	117 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	120 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/call_stmt_1306_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/call_stmt_1306_Sample/crr
      -- CP-element group 118: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/call_stmt_1306_Sample/$entry
      -- 
    crr_2357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(118), ack => call_stmt_1306_call_req_0); -- 
    systemTOP_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(105) & systemTOP_CP_2045_elements(109) & systemTOP_CP_2045_elements(113) & systemTOP_CP_2045_elements(117) & systemTOP_CP_2045_elements(120);
      gj_systemTOP_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	121 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/call_stmt_1306_Update/ccr
      -- CP-element group 119: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/call_stmt_1306_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/call_stmt_1306_update_start_
      -- 
    ccr_2362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(119), ack => call_stmt_1306_call_req_1); -- 
    systemTOP_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= systemTOP_CP_2045_elements(121);
      gj_systemTOP_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: marked-successors 
    -- CP-element group 120: 	103 
    -- CP-element group 120: 	107 
    -- CP-element group 120: 	111 
    -- CP-element group 120: 	115 
    -- CP-element group 120: 	118 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/call_stmt_1306_Sample/cra
      -- CP-element group 120: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/call_stmt_1306_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/call_stmt_1306_sample_completed_
      -- 
    cra_2358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1306_call_ack_0, ack => systemTOP_CP_2045_elements(120)); -- 
    -- CP-element group 121:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	139 
    -- CP-element group 121: marked-successors 
    -- CP-element group 121: 	119 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/call_stmt_1306_Update/cca
      -- CP-element group 121: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/call_stmt_1306_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/call_stmt_1306_update_completed_
      -- 
    cca_2363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1306_call_ack_1, ack => systemTOP_CP_2045_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	86 
    -- CP-element group 122: marked-predecessors 
    -- CP-element group 122: 	124 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1321_Sample/rr
      -- CP-element group 122: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1321_Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1321_sample_start_
      -- 
    rr_2371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(122), ack => type_cast_1321_inst_req_0); -- 
    systemTOP_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(86) & systemTOP_CP_2045_elements(124);
      gj_systemTOP_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	17 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	132 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1321_Update/cr
      -- CP-element group 123: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1321_Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1321_update_start_
      -- 
    cr_2376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(123), ack => type_cast_1321_inst_req_1); -- 
    systemTOP_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(17) & systemTOP_CP_2045_elements(125) & systemTOP_CP_2045_elements(132);
      gj_systemTOP_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: marked-successors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: 	82 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1321_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1321_Sample/ra
      -- CP-element group 124: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1321_sample_completed_
      -- 
    ra_2372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1321_inst_ack_0, ack => systemTOP_CP_2045_elements(124)); -- 
    -- CP-element group 125:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	130 
    -- CP-element group 125: marked-successors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: 	60 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1321_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1321_Update/ca
      -- CP-element group 125: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1321_update_completed_
      -- 
    ca_2377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1321_inst_ack_1, ack => systemTOP_CP_2045_elements(125)); -- 
    -- CP-element group 126:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	65 
    -- CP-element group 126: marked-predecessors 
    -- CP-element group 126: 	128 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1325_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1325_Sample/req
      -- CP-element group 126: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1325_Sample/$entry
      -- 
    req_2385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(126), ack => W_colx_x1x_xi_1307_delayed_1_0_1323_inst_req_0); -- 
    systemTOP_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(65) & systemTOP_CP_2045_elements(128);
      gj_systemTOP_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	17 
    -- CP-element group 127: marked-predecessors 
    -- CP-element group 127: 	129 
    -- CP-element group 127: 	132 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1325_Update/req
      -- CP-element group 127: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1325_update_start_
      -- CP-element group 127: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1325_Update/$entry
      -- 
    req_2390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(127), ack => W_colx_x1x_xi_1307_delayed_1_0_1323_inst_req_1); -- 
    systemTOP_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(17) & systemTOP_CP_2045_elements(129) & systemTOP_CP_2045_elements(132);
      gj_systemTOP_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: marked-successors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: 	61 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1325_sample_completed_
      -- CP-element group 128: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1325_Sample/$exit
      -- CP-element group 128: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1325_Sample/ack
      -- 
    ack_2386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_colx_x1x_xi_1307_delayed_1_0_1323_inst_ack_0, ack => systemTOP_CP_2045_elements(128)); -- 
    -- CP-element group 129:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129: marked-successors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: 	60 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1325_Update/ack
      -- CP-element group 129: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1325_Update/$exit
      -- CP-element group 129: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1325_update_completed_
      -- 
    ack_2391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_colx_x1x_xi_1307_delayed_1_0_1323_inst_ack_1, ack => systemTOP_CP_2045_elements(129)); -- 
    -- CP-element group 130:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	125 
    -- CP-element group 130: 	129 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	132 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1346_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1346_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1346_Sample/rr
      -- 
    rr_2399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(130), ack => type_cast_1346_inst_req_0); -- 
    systemTOP_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(125) & systemTOP_CP_2045_elements(129) & systemTOP_CP_2045_elements(132);
      gj_systemTOP_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	17 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	133 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1346_update_start_
      -- CP-element group 131: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1346_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1346_Update/$entry
      -- 
    cr_2404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(131), ack => type_cast_1346_inst_req_1); -- 
    systemTOP_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(17) & systemTOP_CP_2045_elements(133);
      gj_systemTOP_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: marked-successors 
    -- CP-element group 132: 	123 
    -- CP-element group 132: 	127 
    -- CP-element group 132: 	130 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1346_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1346_Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1346_Sample/ra
      -- 
    ra_2400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1346_inst_ack_0, ack => systemTOP_CP_2045_elements(132)); -- 
    -- CP-element group 133:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	15 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: 	41 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1346_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1346_Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/type_cast_1346_Update/ca
      -- 
    ca_2405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1346_inst_ack_1, ack => systemTOP_CP_2045_elements(133)); -- 
    -- CP-element group 134:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	44 
    -- CP-element group 134: marked-predecessors 
    -- CP-element group 134: 	136 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1350_Sample/req
      -- CP-element group 134: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1350_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1350_sample_start_
      -- 
    req_2413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(134), ack => W_row18x_x1x_xi_1329_delayed_2_0_1348_inst_req_0); -- 
    systemTOP_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(44) & systemTOP_CP_2045_elements(136);
      gj_systemTOP_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 135:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	17 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	137 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1350_Update/req
      -- CP-element group 135: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1350_Update/$entry
      -- CP-element group 135: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1350_update_start_
      -- 
    req_2418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(135), ack => W_row18x_x1x_xi_1329_delayed_2_0_1348_inst_req_1); -- 
    systemTOP_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(17) & systemTOP_CP_2045_elements(137);
      gj_systemTOP_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: marked-successors 
    -- CP-element group 136: 	42 
    -- CP-element group 136: 	134 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1350_Sample/ack
      -- CP-element group 136: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1350_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1350_sample_completed_
      -- 
    ack_2414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_row18x_x1x_xi_1329_delayed_2_0_1348_inst_ack_0, ack => systemTOP_CP_2045_elements(136)); -- 
    -- CP-element group 137:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	15 
    -- CP-element group 137: marked-successors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: 	41 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1350_Update/ack
      -- CP-element group 137: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1350_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/assign_stmt_1350_update_completed_
      -- 
    ack_2419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_row18x_x1x_xi_1329_delayed_2_0_1348_inst_ack_1, ack => systemTOP_CP_2045_elements(137)); -- 
    -- CP-element group 138:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	14 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	15 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group systemTOP_CP_2045_elements(138) is a control-delay.
    cp_element_138_delay: control_delay_element  generic map(name => " 138_delay", delay_value => 1)  port map(req => systemTOP_CP_2045_elements(14), ack => systemTOP_CP_2045_elements(138), clk => clk, reset =>reset);
    -- CP-element group 139:  join  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	121 
    -- CP-element group 139: 	17 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	11 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_1191/do_while_stmt_1218/do_while_stmt_1218_loop_body/$exit
      -- 
    systemTOP_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(121) & systemTOP_CP_2045_elements(17);
      gj_systemTOP_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	10 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (2) 
      -- CP-element group 140: 	 branch_block_stmt_1191/do_while_stmt_1218/loop_exit/ack
      -- CP-element group 140: 	 branch_block_stmt_1191/do_while_stmt_1218/loop_exit/$exit
      -- 
    ack_2424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1218_branch_ack_0, ack => systemTOP_CP_2045_elements(140)); -- 
    -- CP-element group 141:  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	10 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (2) 
      -- CP-element group 141: 	 branch_block_stmt_1191/do_while_stmt_1218/loop_taken/ack
      -- CP-element group 141: 	 branch_block_stmt_1191/do_while_stmt_1218/loop_taken/$exit
      -- 
    ack_2428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1218_branch_ack_1, ack => systemTOP_CP_2045_elements(141)); -- 
    -- CP-element group 142:  transition  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	8 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	1 
    -- CP-element group 142:  members (1) 
      -- CP-element group 142: 	 branch_block_stmt_1191/do_while_stmt_1218/$exit
      -- 
    systemTOP_CP_2045_elements(142) <= systemTOP_CP_2045_elements(8);
    -- CP-element group 143:  fork  transition  place  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	1 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	205 
    -- CP-element group 143: 	206 
    -- CP-element group 143:  members (12) 
      -- CP-element group 143: 	 branch_block_stmt_1191/whilex_xbodyx_xi_maxPool3Dx_xexit
      -- CP-element group 143: 	 branch_block_stmt_1191/if_stmt_1381_if_link/if_choice_transition
      -- CP-element group 143: 	 branch_block_stmt_1191/if_stmt_1381_if_link/$exit
      -- CP-element group 143: 	 branch_block_stmt_1191/whilex_xbodyx_xi_maxPool3Dx_xexit_PhiReq/$entry
      -- CP-element group 143: 	 branch_block_stmt_1191/whilex_xbodyx_xi_maxPool3Dx_xexit_PhiReq/phi_stmt_1386/$entry
      -- CP-element group 143: 	 branch_block_stmt_1191/whilex_xbodyx_xi_maxPool3Dx_xexit_PhiReq/phi_stmt_1386/phi_stmt_1386_sources/$entry
      -- CP-element group 143: 	 branch_block_stmt_1191/whilex_xbodyx_xi_maxPool3Dx_xexit_PhiReq/phi_stmt_1386/phi_stmt_1386_sources/type_cast_1389/$entry
      -- CP-element group 143: 	 branch_block_stmt_1191/whilex_xbodyx_xi_maxPool3Dx_xexit_PhiReq/phi_stmt_1386/phi_stmt_1386_sources/type_cast_1389/SplitProtocol/$entry
      -- CP-element group 143: 	 branch_block_stmt_1191/whilex_xbodyx_xi_maxPool3Dx_xexit_PhiReq/phi_stmt_1386/phi_stmt_1386_sources/type_cast_1389/SplitProtocol/Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_1191/whilex_xbodyx_xi_maxPool3Dx_xexit_PhiReq/phi_stmt_1386/phi_stmt_1386_sources/type_cast_1389/SplitProtocol/Sample/rr
      -- CP-element group 143: 	 branch_block_stmt_1191/whilex_xbodyx_xi_maxPool3Dx_xexit_PhiReq/phi_stmt_1386/phi_stmt_1386_sources/type_cast_1389/SplitProtocol/Update/$entry
      -- CP-element group 143: 	 branch_block_stmt_1191/whilex_xbodyx_xi_maxPool3Dx_xexit_PhiReq/phi_stmt_1386/phi_stmt_1386_sources/type_cast_1389/SplitProtocol/Update/cr
      -- 
    if_choice_transition_2442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1381_branch_ack_1, ack => systemTOP_CP_2045_elements(143)); -- 
    rr_2788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(143), ack => type_cast_1389_inst_req_0); -- 
    cr_2793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(143), ack => type_cast_1389_inst_req_1); -- 
    -- CP-element group 144:  merge  transition  place  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	1 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (5) 
      -- CP-element group 144: 	 branch_block_stmt_1191/if_stmt_1381_else_link/else_choice_transition
      -- CP-element group 144: 	 branch_block_stmt_1191/if_stmt_1381_else_link/$exit
      -- CP-element group 144: 	 branch_block_stmt_1191/if_stmt_1381__exit__
      -- CP-element group 144: 	 branch_block_stmt_1191/merge_stmt_1385__entry__
      -- CP-element group 144: 	 branch_block_stmt_1191/merge_stmt_1385_dead_link/$entry
      -- 
    else_choice_transition_2446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1381_branch_ack_0, ack => systemTOP_CP_2045_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	208 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1395_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1395_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1395_sample_completed_
      -- 
    ra_2459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1395_inst_ack_0, ack => systemTOP_CP_2045_elements(145)); -- 
    -- CP-element group 146:  fork  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	208 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	155 
    -- CP-element group 146: 	158 
    -- CP-element group 146: 	161 
    -- CP-element group 146: 	164 
    -- CP-element group 146: 	167 
    -- CP-element group 146: 	170 
    -- CP-element group 146: 	173 
    -- CP-element group 146: 	176 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1395_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1395_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1395_Update/$exit
      -- 
    ca_2464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1395_inst_ack_1, ack => systemTOP_CP_2045_elements(146)); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	208 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1399_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1399_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1399_sample_completed_
      -- 
    ra_2473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1399_inst_ack_0, ack => systemTOP_CP_2045_elements(147)); -- 
    -- CP-element group 148:  transition  input  output  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	208 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	149 
    -- CP-element group 148:  members (6) 
      -- CP-element group 148: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1399_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1399_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1399_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1401_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1401_Sample/$entry
      -- CP-element group 148: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1401_Sample/req
      -- 
    ca_2478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1399_inst_ack_1, ack => systemTOP_CP_2045_elements(148)); -- 
    req_2486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(148), ack => WPIPE_system_output_pipe_1401_inst_req_0); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	148 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1401_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1401_update_start_
      -- CP-element group 149: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1401_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1401_Sample/ack
      -- CP-element group 149: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1401_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1401_Update/req
      -- 
    ack_2487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1401_inst_ack_0, ack => systemTOP_CP_2045_elements(149)); -- 
    req_2491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(149), ack => WPIPE_system_output_pipe_1401_inst_req_1); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	179 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1401_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1401_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1401_Update/ack
      -- 
    ack_2492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1401_inst_ack_1, ack => systemTOP_CP_2045_elements(150)); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	208 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1405_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1405_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1405_Sample/cra
      -- 
    cra_2501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1405_call_ack_0, ack => systemTOP_CP_2045_elements(151)); -- 
    -- CP-element group 152:  transition  input  output  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	208 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152:  members (6) 
      -- CP-element group 152: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1405_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1405_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1405_Update/cca
      -- CP-element group 152: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1409_sample_start_
      -- CP-element group 152: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1409_Sample/$entry
      -- CP-element group 152: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1409_Sample/rr
      -- 
    cca_2506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1405_call_ack_1, ack => systemTOP_CP_2045_elements(152)); -- 
    rr_2514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(152), ack => type_cast_1409_inst_req_0); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	152 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1409_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1409_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1409_Sample/ra
      -- 
    ra_2515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1409_inst_ack_0, ack => systemTOP_CP_2045_elements(153)); -- 
    -- CP-element group 154:  fork  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	208 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154: 	158 
    -- CP-element group 154: 	161 
    -- CP-element group 154: 	164 
    -- CP-element group 154: 	167 
    -- CP-element group 154: 	170 
    -- CP-element group 154: 	173 
    -- CP-element group 154: 	176 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1409_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1409_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1409_Update/ca
      -- 
    ca_2520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1409_inst_ack_1, ack => systemTOP_CP_2045_elements(154)); -- 
    -- CP-element group 155:  join  transition  output  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: 	146 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1418_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1418_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1418_Sample/rr
      -- 
    rr_2528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(155), ack => type_cast_1418_inst_req_0); -- 
    systemTOP_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(154) & systemTOP_CP_2045_elements(146);
      gj_systemTOP_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1418_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1418_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1418_Sample/ra
      -- 
    ra_2529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1418_inst_ack_0, ack => systemTOP_CP_2045_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	208 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	200 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1418_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1418_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1418_Update/ca
      -- 
    ca_2534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1418_inst_ack_1, ack => systemTOP_CP_2045_elements(157)); -- 
    -- CP-element group 158:  join  transition  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	154 
    -- CP-element group 158: 	146 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1428_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1428_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1428_Sample/rr
      -- 
    rr_2542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(158), ack => type_cast_1428_inst_req_0); -- 
    systemTOP_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(154) & systemTOP_CP_2045_elements(146);
      gj_systemTOP_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1428_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1428_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1428_Sample/ra
      -- 
    ra_2543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1428_inst_ack_0, ack => systemTOP_CP_2045_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	208 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	197 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1428_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1428_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1428_Update/ca
      -- 
    ca_2548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1428_inst_ack_1, ack => systemTOP_CP_2045_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	154 
    -- CP-element group 161: 	146 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1438_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1438_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1438_Sample/rr
      -- 
    rr_2556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(161), ack => type_cast_1438_inst_req_0); -- 
    systemTOP_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(154) & systemTOP_CP_2045_elements(146);
      gj_systemTOP_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1438_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1438_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1438_Sample/ra
      -- 
    ra_2557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1438_inst_ack_0, ack => systemTOP_CP_2045_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	208 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	194 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1438_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1438_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1438_Update/ca
      -- 
    ca_2562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1438_inst_ack_1, ack => systemTOP_CP_2045_elements(163)); -- 
    -- CP-element group 164:  join  transition  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	154 
    -- CP-element group 164: 	146 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1448_sample_start_
      -- CP-element group 164: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1448_Sample/$entry
      -- CP-element group 164: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1448_Sample/rr
      -- 
    rr_2570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(164), ack => type_cast_1448_inst_req_0); -- 
    systemTOP_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(154) & systemTOP_CP_2045_elements(146);
      gj_systemTOP_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1448_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1448_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1448_Sample/ra
      -- 
    ra_2571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1448_inst_ack_0, ack => systemTOP_CP_2045_elements(165)); -- 
    -- CP-element group 166:  transition  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	208 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	191 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1448_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1448_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1448_Update/ca
      -- 
    ca_2576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1448_inst_ack_1, ack => systemTOP_CP_2045_elements(166)); -- 
    -- CP-element group 167:  join  transition  output  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	154 
    -- CP-element group 167: 	146 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	168 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1458_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1458_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1458_Sample/rr
      -- 
    rr_2584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(167), ack => type_cast_1458_inst_req_0); -- 
    systemTOP_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(154) & systemTOP_CP_2045_elements(146);
      gj_systemTOP_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	167 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1458_sample_completed_
      -- CP-element group 168: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1458_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1458_Sample/ra
      -- 
    ra_2585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1458_inst_ack_0, ack => systemTOP_CP_2045_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	208 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	188 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1458_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1458_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1458_Update/ca
      -- 
    ca_2590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1458_inst_ack_1, ack => systemTOP_CP_2045_elements(169)); -- 
    -- CP-element group 170:  join  transition  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	154 
    -- CP-element group 170: 	146 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1468_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1468_Sample/$entry
      -- CP-element group 170: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1468_Sample/rr
      -- 
    rr_2598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(170), ack => type_cast_1468_inst_req_0); -- 
    systemTOP_cp_element_group_170: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_170"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(154) & systemTOP_CP_2045_elements(146);
      gj_systemTOP_cp_element_group_170 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(170), clk => clk, reset => reset); --
    end block;
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1468_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1468_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1468_Sample/ra
      -- 
    ra_2599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1468_inst_ack_0, ack => systemTOP_CP_2045_elements(171)); -- 
    -- CP-element group 172:  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	208 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	185 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1468_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1468_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1468_Update/ca
      -- 
    ca_2604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1468_inst_ack_1, ack => systemTOP_CP_2045_elements(172)); -- 
    -- CP-element group 173:  join  transition  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	154 
    -- CP-element group 173: 	146 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1478_sample_start_
      -- CP-element group 173: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1478_Sample/$entry
      -- CP-element group 173: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1478_Sample/rr
      -- 
    rr_2612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(173), ack => type_cast_1478_inst_req_0); -- 
    systemTOP_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(154) & systemTOP_CP_2045_elements(146);
      gj_systemTOP_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1478_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1478_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1478_Sample/ra
      -- 
    ra_2613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1478_inst_ack_0, ack => systemTOP_CP_2045_elements(174)); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	208 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	182 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1478_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1478_Update/$exit
      -- CP-element group 175: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1478_Update/ca
      -- 
    ca_2618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1478_inst_ack_1, ack => systemTOP_CP_2045_elements(175)); -- 
    -- CP-element group 176:  join  transition  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	154 
    -- CP-element group 176: 	146 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1488_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1488_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1488_Sample/rr
      -- 
    rr_2626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(176), ack => type_cast_1488_inst_req_0); -- 
    systemTOP_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(154) & systemTOP_CP_2045_elements(146);
      gj_systemTOP_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1488_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1488_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1488_Sample/ra
      -- 
    ra_2627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1488_inst_ack_0, ack => systemTOP_CP_2045_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	208 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1488_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1488_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1488_Update/ca
      -- 
    ca_2632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1488_inst_ack_1, ack => systemTOP_CP_2045_elements(178)); -- 
    -- CP-element group 179:  join  transition  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: 	150 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1490_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1490_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1490_Sample/req
      -- 
    req_2640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(179), ack => WPIPE_system_output_pipe_1490_inst_req_0); -- 
    systemTOP_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(178) & systemTOP_CP_2045_elements(150);
      gj_systemTOP_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (6) 
      -- CP-element group 180: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1490_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1490_update_start_
      -- CP-element group 180: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1490_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1490_Sample/ack
      -- CP-element group 180: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1490_Update/$entry
      -- CP-element group 180: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1490_Update/req
      -- 
    ack_2641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1490_inst_ack_0, ack => systemTOP_CP_2045_elements(180)); -- 
    req_2645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(180), ack => WPIPE_system_output_pipe_1490_inst_req_1); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1490_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1490_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1490_Update/ack
      -- 
    ack_2646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1490_inst_ack_1, ack => systemTOP_CP_2045_elements(181)); -- 
    -- CP-element group 182:  join  transition  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	175 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1493_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1493_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1493_Sample/req
      -- 
    req_2654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(182), ack => WPIPE_system_output_pipe_1493_inst_req_0); -- 
    systemTOP_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(175) & systemTOP_CP_2045_elements(181);
      gj_systemTOP_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  transition  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183:  members (6) 
      -- CP-element group 183: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1493_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1493_update_start_
      -- CP-element group 183: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1493_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1493_Sample/ack
      -- CP-element group 183: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1493_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1493_Update/req
      -- 
    ack_2655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1493_inst_ack_0, ack => systemTOP_CP_2045_elements(183)); -- 
    req_2659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(183), ack => WPIPE_system_output_pipe_1493_inst_req_1); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1493_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1493_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1493_Update/ack
      -- 
    ack_2660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1493_inst_ack_1, ack => systemTOP_CP_2045_elements(184)); -- 
    -- CP-element group 185:  join  transition  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	172 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1496_sample_start_
      -- CP-element group 185: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1496_Sample/$entry
      -- CP-element group 185: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1496_Sample/req
      -- 
    req_2668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(185), ack => WPIPE_system_output_pipe_1496_inst_req_0); -- 
    systemTOP_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(172) & systemTOP_CP_2045_elements(184);
      gj_systemTOP_cp_element_group_185 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (6) 
      -- CP-element group 186: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1496_sample_completed_
      -- CP-element group 186: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1496_update_start_
      -- CP-element group 186: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1496_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1496_Sample/ack
      -- CP-element group 186: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1496_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1496_Update/req
      -- 
    ack_2669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1496_inst_ack_0, ack => systemTOP_CP_2045_elements(186)); -- 
    req_2673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(186), ack => WPIPE_system_output_pipe_1496_inst_req_1); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1496_update_completed_
      -- CP-element group 187: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1496_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1496_Update/ack
      -- 
    ack_2674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1496_inst_ack_1, ack => systemTOP_CP_2045_elements(187)); -- 
    -- CP-element group 188:  join  transition  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	169 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1499_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1499_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1499_Sample/req
      -- 
    req_2682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(188), ack => WPIPE_system_output_pipe_1499_inst_req_0); -- 
    systemTOP_cp_element_group_188: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_188"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(169) & systemTOP_CP_2045_elements(187);
      gj_systemTOP_cp_element_group_188 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(188), clk => clk, reset => reset); --
    end block;
    -- CP-element group 189:  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (6) 
      -- CP-element group 189: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1499_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1499_update_start_
      -- CP-element group 189: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1499_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1499_Sample/ack
      -- CP-element group 189: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1499_Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1499_Update/req
      -- 
    ack_2683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1499_inst_ack_0, ack => systemTOP_CP_2045_elements(189)); -- 
    req_2687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(189), ack => WPIPE_system_output_pipe_1499_inst_req_1); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1499_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1499_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1499_Update/ack
      -- 
    ack_2688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1499_inst_ack_1, ack => systemTOP_CP_2045_elements(190)); -- 
    -- CP-element group 191:  join  transition  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	166 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1502_sample_start_
      -- CP-element group 191: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1502_Sample/$entry
      -- CP-element group 191: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1502_Sample/req
      -- 
    req_2696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(191), ack => WPIPE_system_output_pipe_1502_inst_req_0); -- 
    systemTOP_cp_element_group_191: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_191"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(166) & systemTOP_CP_2045_elements(190);
      gj_systemTOP_cp_element_group_191 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(191), clk => clk, reset => reset); --
    end block;
    -- CP-element group 192:  transition  input  output  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192:  members (6) 
      -- CP-element group 192: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1502_sample_completed_
      -- CP-element group 192: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1502_update_start_
      -- CP-element group 192: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1502_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1502_Sample/ack
      -- CP-element group 192: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1502_Update/$entry
      -- CP-element group 192: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1502_Update/req
      -- 
    ack_2697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1502_inst_ack_0, ack => systemTOP_CP_2045_elements(192)); -- 
    req_2701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(192), ack => WPIPE_system_output_pipe_1502_inst_req_1); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1502_update_completed_
      -- CP-element group 193: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1502_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1502_Update/ack
      -- 
    ack_2702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1502_inst_ack_1, ack => systemTOP_CP_2045_elements(193)); -- 
    -- CP-element group 194:  join  transition  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	163 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1505_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1505_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1505_Sample/req
      -- 
    req_2710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(194), ack => WPIPE_system_output_pipe_1505_inst_req_0); -- 
    systemTOP_cp_element_group_194: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_194"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(163) & systemTOP_CP_2045_elements(193);
      gj_systemTOP_cp_element_group_194 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(194), clk => clk, reset => reset); --
    end block;
    -- CP-element group 195:  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (6) 
      -- CP-element group 195: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1505_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1505_update_start_
      -- CP-element group 195: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1505_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1505_Sample/ack
      -- CP-element group 195: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1505_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1505_Update/req
      -- 
    ack_2711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1505_inst_ack_0, ack => systemTOP_CP_2045_elements(195)); -- 
    req_2715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(195), ack => WPIPE_system_output_pipe_1505_inst_req_1); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	197 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1505_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1505_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1505_Update/ack
      -- 
    ack_2716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1505_inst_ack_1, ack => systemTOP_CP_2045_elements(196)); -- 
    -- CP-element group 197:  join  transition  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	160 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1508_sample_start_
      -- CP-element group 197: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1508_Sample/$entry
      -- CP-element group 197: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1508_Sample/req
      -- 
    req_2724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(197), ack => WPIPE_system_output_pipe_1508_inst_req_0); -- 
    systemTOP_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(160) & systemTOP_CP_2045_elements(196);
      gj_systemTOP_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198:  members (6) 
      -- CP-element group 198: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1508_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1508_update_start_
      -- CP-element group 198: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1508_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1508_Sample/ack
      -- CP-element group 198: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1508_Update/$entry
      -- CP-element group 198: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1508_Update/req
      -- 
    ack_2725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1508_inst_ack_0, ack => systemTOP_CP_2045_elements(198)); -- 
    req_2729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(198), ack => WPIPE_system_output_pipe_1508_inst_req_1); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1508_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1508_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1508_Update/ack
      -- 
    ack_2730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1508_inst_ack_1, ack => systemTOP_CP_2045_elements(199)); -- 
    -- CP-element group 200:  join  transition  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	157 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1511_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1511_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1511_Sample/req
      -- 
    req_2738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(200), ack => WPIPE_system_output_pipe_1511_inst_req_0); -- 
    systemTOP_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(157) & systemTOP_CP_2045_elements(199);
      gj_systemTOP_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1511_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1511_update_start_
      -- CP-element group 201: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1511_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1511_Sample/ack
      -- CP-element group 201: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1511_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1511_Update/req
      -- 
    ack_2739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1511_inst_ack_0, ack => systemTOP_CP_2045_elements(201)); -- 
    req_2743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(201), ack => WPIPE_system_output_pipe_1511_inst_req_1); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1511_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1511_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/WPIPE_system_output_pipe_1511_Update/ack
      -- CP-element group 202: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1514_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1514_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1514_Sample/crr
      -- 
    ack_2744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_system_output_pipe_1511_inst_ack_1, ack => systemTOP_CP_2045_elements(202)); -- 
    crr_2752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(202), ack => call_stmt_1514_call_req_0); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1514_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1514_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1514_Sample/cra
      -- 
    cra_2753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1514_call_ack_0, ack => systemTOP_CP_2045_elements(203)); -- 
    -- CP-element group 204:  transition  place  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	208 
    -- CP-element group 204: successors 
    -- CP-element group 204:  members (16) 
      -- CP-element group 204: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/$exit
      -- CP-element group 204: 	 $exit
      -- CP-element group 204: 	 branch_block_stmt_1191/$exit
      -- CP-element group 204: 	 branch_block_stmt_1191/branch_block_stmt_1191__exit__
      -- CP-element group 204: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514__exit__
      -- CP-element group 204: 	 branch_block_stmt_1191/return__
      -- CP-element group 204: 	 branch_block_stmt_1191/merge_stmt_1516__exit__
      -- CP-element group 204: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1514_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1514_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1514_Update/cca
      -- CP-element group 204: 	 branch_block_stmt_1191/return___PhiReq/$entry
      -- CP-element group 204: 	 branch_block_stmt_1191/return___PhiReq/$exit
      -- CP-element group 204: 	 branch_block_stmt_1191/merge_stmt_1516_PhiReqMerge
      -- CP-element group 204: 	 branch_block_stmt_1191/merge_stmt_1516_PhiAck/$entry
      -- CP-element group 204: 	 branch_block_stmt_1191/merge_stmt_1516_PhiAck/$exit
      -- CP-element group 204: 	 branch_block_stmt_1191/merge_stmt_1516_PhiAck/dummy
      -- 
    cca_2758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1514_call_ack_1, ack => systemTOP_CP_2045_elements(204)); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	143 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	207 
    -- CP-element group 205:  members (2) 
      -- CP-element group 205: 	 branch_block_stmt_1191/whilex_xbodyx_xi_maxPool3Dx_xexit_PhiReq/phi_stmt_1386/phi_stmt_1386_sources/type_cast_1389/SplitProtocol/Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_1191/whilex_xbodyx_xi_maxPool3Dx_xexit_PhiReq/phi_stmt_1386/phi_stmt_1386_sources/type_cast_1389/SplitProtocol/Sample/ra
      -- 
    ra_2789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1389_inst_ack_0, ack => systemTOP_CP_2045_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	143 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (2) 
      -- CP-element group 206: 	 branch_block_stmt_1191/whilex_xbodyx_xi_maxPool3Dx_xexit_PhiReq/phi_stmt_1386/phi_stmt_1386_sources/type_cast_1389/SplitProtocol/Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_1191/whilex_xbodyx_xi_maxPool3Dx_xexit_PhiReq/phi_stmt_1386/phi_stmt_1386_sources/type_cast_1389/SplitProtocol/Update/ca
      -- 
    ca_2794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1389_inst_ack_1, ack => systemTOP_CP_2045_elements(206)); -- 
    -- CP-element group 207:  join  transition  place  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	205 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (8) 
      -- CP-element group 207: 	 branch_block_stmt_1191/whilex_xbodyx_xi_maxPool3Dx_xexit_PhiReq/$exit
      -- CP-element group 207: 	 branch_block_stmt_1191/whilex_xbodyx_xi_maxPool3Dx_xexit_PhiReq/phi_stmt_1386/$exit
      -- CP-element group 207: 	 branch_block_stmt_1191/whilex_xbodyx_xi_maxPool3Dx_xexit_PhiReq/phi_stmt_1386/phi_stmt_1386_sources/$exit
      -- CP-element group 207: 	 branch_block_stmt_1191/whilex_xbodyx_xi_maxPool3Dx_xexit_PhiReq/phi_stmt_1386/phi_stmt_1386_sources/type_cast_1389/$exit
      -- CP-element group 207: 	 branch_block_stmt_1191/whilex_xbodyx_xi_maxPool3Dx_xexit_PhiReq/phi_stmt_1386/phi_stmt_1386_sources/type_cast_1389/SplitProtocol/$exit
      -- CP-element group 207: 	 branch_block_stmt_1191/whilex_xbodyx_xi_maxPool3Dx_xexit_PhiReq/phi_stmt_1386/phi_stmt_1386_req
      -- CP-element group 207: 	 branch_block_stmt_1191/merge_stmt_1385_PhiReqMerge
      -- CP-element group 207: 	 branch_block_stmt_1191/merge_stmt_1385_PhiAck/$entry
      -- 
    phi_stmt_1386_req_2795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1386_req_2795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(207), ack => phi_stmt_1386_req_0); -- 
    systemTOP_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "systemTOP_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= systemTOP_CP_2045_elements(205) & systemTOP_CP_2045_elements(206);
      gj_systemTOP_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => systemTOP_CP_2045_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	152 
    -- CP-element group 208: 	154 
    -- CP-element group 208: 	157 
    -- CP-element group 208: 	160 
    -- CP-element group 208: 	163 
    -- CP-element group 208: 	166 
    -- CP-element group 208: 	169 
    -- CP-element group 208: 	172 
    -- CP-element group 208: 	175 
    -- CP-element group 208: 	178 
    -- CP-element group 208: 	145 
    -- CP-element group 208: 	146 
    -- CP-element group 208: 	147 
    -- CP-element group 208: 	148 
    -- CP-element group 208: 	151 
    -- CP-element group 208: 	204 
    -- CP-element group 208:  members (53) 
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1399_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1399_Sample/rr
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1399_Sample/$entry
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1399_Update/cr
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1399_update_start_
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1395_Sample/rr
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1395_Sample/$entry
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1395_update_start_
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1395_sample_start_
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/$entry
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1399_sample_start_
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1395_Update/cr
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1395_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_1191/merge_stmt_1385__exit__
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514__entry__
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1405_sample_start_
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1405_update_start_
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1405_Sample/$entry
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1405_Sample/crr
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1405_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1405_Update/ccr
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1409_update_start_
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1409_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1409_Update/cr
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1418_update_start_
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1418_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1418_Update/cr
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1428_update_start_
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1428_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1428_Update/cr
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1438_update_start_
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1438_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1438_Update/cr
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1448_update_start_
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1448_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1448_Update/cr
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1458_update_start_
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1458_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1458_Update/cr
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1468_update_start_
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1468_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1468_Update/cr
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1478_update_start_
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1478_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1478_Update/cr
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1488_update_start_
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1488_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/type_cast_1488_Update/cr
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1514_update_start_
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1514_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_1191/assign_stmt_1396_to_call_stmt_1514/call_stmt_1514_Update/ccr
      -- CP-element group 208: 	 branch_block_stmt_1191/merge_stmt_1385_PhiAck/$exit
      -- CP-element group 208: 	 branch_block_stmt_1191/merge_stmt_1385_PhiAck/phi_stmt_1386_ack
      -- 
    phi_stmt_1386_ack_2800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1386_ack_0, ack => systemTOP_CP_2045_elements(208)); -- 
    rr_2472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(208), ack => type_cast_1399_inst_req_0); -- 
    cr_2477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(208), ack => type_cast_1399_inst_req_1); -- 
    rr_2458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(208), ack => type_cast_1395_inst_req_0); -- 
    cr_2463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(208), ack => type_cast_1395_inst_req_1); -- 
    crr_2500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(208), ack => call_stmt_1405_call_req_0); -- 
    ccr_2505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(208), ack => call_stmt_1405_call_req_1); -- 
    cr_2519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(208), ack => type_cast_1409_inst_req_1); -- 
    cr_2533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(208), ack => type_cast_1418_inst_req_1); -- 
    cr_2547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(208), ack => type_cast_1428_inst_req_1); -- 
    cr_2561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(208), ack => type_cast_1438_inst_req_1); -- 
    cr_2575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(208), ack => type_cast_1448_inst_req_1); -- 
    cr_2589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(208), ack => type_cast_1458_inst_req_1); -- 
    cr_2603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(208), ack => type_cast_1468_inst_req_1); -- 
    cr_2617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(208), ack => type_cast_1478_inst_req_1); -- 
    cr_2631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(208), ack => type_cast_1488_inst_req_1); -- 
    ccr_2757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => systemTOP_CP_2045_elements(208), ack => call_stmt_1514_call_req_1); -- 
    systemTOP_do_while_stmt_1218_terminator_2429: loop_terminator -- 
      generic map (name => " systemTOP_do_while_stmt_1218_terminator_2429", max_iterations_in_flight =>15) 
      port map(loop_body_exit => systemTOP_CP_2045_elements(11),loop_continue => systemTOP_CP_2045_elements(141),loop_terminate => systemTOP_CP_2045_elements(140),loop_back => systemTOP_CP_2045_elements(9),loop_exit => systemTOP_CP_2045_elements(8),clk => clk, reset => reset); -- 
    phi_stmt_1220_phi_seq_2161_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= systemTOP_CP_2045_elements(26);
      systemTOP_CP_2045_elements(31)<= src_sample_reqs(0);
      src_sample_acks(0)  <= systemTOP_CP_2045_elements(35);
      systemTOP_CP_2045_elements(32)<= src_update_reqs(0);
      src_update_acks(0)  <= systemTOP_CP_2045_elements(36);
      systemTOP_CP_2045_elements(27) <= phi_mux_reqs(0);
      triggers(1)  <= systemTOP_CP_2045_elements(28);
      systemTOP_CP_2045_elements(37)<= src_sample_reqs(1);
      src_sample_acks(1)  <= systemTOP_CP_2045_elements(37);
      systemTOP_CP_2045_elements(38)<= src_update_reqs(1);
      src_update_acks(1)  <= systemTOP_CP_2045_elements(39);
      systemTOP_CP_2045_elements(29) <= phi_mux_reqs(1);
      phi_stmt_1220_phi_seq_2161 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1220_phi_seq_2161") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => systemTOP_CP_2045_elements(22), 
          phi_sample_ack => systemTOP_CP_2045_elements(23), 
          phi_update_req => systemTOP_CP_2045_elements(24), 
          phi_update_ack => systemTOP_CP_2045_elements(25), 
          phi_mux_ack => systemTOP_CP_2045_elements(30), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1225_phi_seq_2205_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= systemTOP_CP_2045_elements(45);
      systemTOP_CP_2045_elements(50)<= src_sample_reqs(0);
      src_sample_acks(0)  <= systemTOP_CP_2045_elements(54);
      systemTOP_CP_2045_elements(51)<= src_update_reqs(0);
      src_update_acks(0)  <= systemTOP_CP_2045_elements(55);
      systemTOP_CP_2045_elements(46) <= phi_mux_reqs(0);
      triggers(1)  <= systemTOP_CP_2045_elements(47);
      systemTOP_CP_2045_elements(56)<= src_sample_reqs(1);
      src_sample_acks(1)  <= systemTOP_CP_2045_elements(56);
      systemTOP_CP_2045_elements(57)<= src_update_reqs(1);
      src_update_acks(1)  <= systemTOP_CP_2045_elements(58);
      systemTOP_CP_2045_elements(48) <= phi_mux_reqs(1);
      phi_stmt_1225_phi_seq_2205 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1225_phi_seq_2205") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => systemTOP_CP_2045_elements(16), 
          phi_sample_ack => systemTOP_CP_2045_elements(43), 
          phi_update_req => systemTOP_CP_2045_elements(18), 
          phi_update_ack => systemTOP_CP_2045_elements(44), 
          phi_mux_ack => systemTOP_CP_2045_elements(49), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1230_phi_seq_2249_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= systemTOP_CP_2045_elements(66);
      systemTOP_CP_2045_elements(71)<= src_sample_reqs(0);
      src_sample_acks(0)  <= systemTOP_CP_2045_elements(75);
      systemTOP_CP_2045_elements(72)<= src_update_reqs(0);
      src_update_acks(0)  <= systemTOP_CP_2045_elements(76);
      systemTOP_CP_2045_elements(67) <= phi_mux_reqs(0);
      triggers(1)  <= systemTOP_CP_2045_elements(68);
      systemTOP_CP_2045_elements(77)<= src_sample_reqs(1);
      src_sample_acks(1)  <= systemTOP_CP_2045_elements(77);
      systemTOP_CP_2045_elements(78)<= src_update_reqs(1);
      src_update_acks(1)  <= systemTOP_CP_2045_elements(79);
      systemTOP_CP_2045_elements(69) <= phi_mux_reqs(1);
      phi_stmt_1230_phi_seq_2249 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1230_phi_seq_2249") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => systemTOP_CP_2045_elements(62), 
          phi_sample_ack => systemTOP_CP_2045_elements(63), 
          phi_update_req => systemTOP_CP_2045_elements(64), 
          phi_update_ack => systemTOP_CP_2045_elements(65), 
          phi_mux_ack => systemTOP_CP_2045_elements(70), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1235_phi_seq_2293_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= systemTOP_CP_2045_elements(87);
      systemTOP_CP_2045_elements(92)<= src_sample_reqs(0);
      src_sample_acks(0)  <= systemTOP_CP_2045_elements(96);
      systemTOP_CP_2045_elements(93)<= src_update_reqs(0);
      src_update_acks(0)  <= systemTOP_CP_2045_elements(97);
      systemTOP_CP_2045_elements(88) <= phi_mux_reqs(0);
      triggers(1)  <= systemTOP_CP_2045_elements(89);
      systemTOP_CP_2045_elements(98)<= src_sample_reqs(1);
      src_sample_acks(1)  <= systemTOP_CP_2045_elements(98);
      systemTOP_CP_2045_elements(99)<= src_update_reqs(1);
      src_update_acks(1)  <= systemTOP_CP_2045_elements(100);
      systemTOP_CP_2045_elements(90) <= phi_mux_reqs(1);
      phi_stmt_1235_phi_seq_2293 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1235_phi_seq_2293") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => systemTOP_CP_2045_elements(83), 
          phi_sample_ack => systemTOP_CP_2045_elements(84), 
          phi_update_req => systemTOP_CP_2045_elements(85), 
          phi_update_ack => systemTOP_CP_2045_elements(86), 
          phi_mux_ack => systemTOP_CP_2045_elements(91), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2113_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= systemTOP_CP_2045_elements(12);
        preds(1)  <= systemTOP_CP_2045_elements(13);
        entry_tmerge_2113 : transition_merge -- 
          generic map(name => " entry_tmerge_2113")
          port map (preds => preds, symbol_out => systemTOP_CP_2045_elements(14));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal NOT_u1_u1_1380_wire : std_logic_vector(0 downto 0);
    signal add41x_xi_1263 : std_logic_vector(31 downto 0);
    signal add43x_xi_1274 : std_logic_vector(31 downto 0);
    signal add50x_xi_1280 : std_logic_vector(31 downto 0);
    signal add54x_xi_1286 : std_logic_vector(31 downto 0);
    signal add57x_xi_1292 : std_logic_vector(31 downto 0);
    signal add79x_xi_1368 : std_logic_vector(31 downto 0);
    signal call1_1405 : std_logic_vector(63 downto 0);
    signal call_1194 : std_logic_vector(63 downto 0);
    signal callx_xi_1306 : std_logic_vector(7 downto 0);
    signal chlx_x0x_xi_1235 : std_logic_vector(15 downto 0);
    signal chlx_x0x_xi_at_entry_1212 : std_logic_vector(15 downto 0);
    signal chlx_x1x_xi_1337 : std_logic_vector(15 downto 0);
    signal cmp72x_xi_1343 : std_logic_vector(0 downto 0);
    signal cmp84x_xi_1374 : std_logic_vector(0 downto 0);
    signal cmpx_xi_1318 : std_logic_vector(0 downto 0);
    signal colx_x1x_xi_1230 : std_logic_vector(15 downto 0);
    signal colx_x1x_xi_1307_delayed_1_0_1325 : std_logic_vector(15 downto 0);
    signal colx_x1x_xi_at_entry_1207 : std_logic_vector(15 downto 0);
    signal colx_x2x_xi_1362 : std_logic_vector(15 downto 0);
    signal conv10_1429 : std_logic_vector(7 downto 0);
    signal conv16_1439 : std_logic_vector(7 downto 0);
    signal conv22_1449 : std_logic_vector(7 downto 0);
    signal conv28_1459 : std_logic_vector(7 downto 0);
    signal conv2_1410 : std_logic_vector(63 downto 0);
    signal conv31x_xi_1244 : std_logic_vector(31 downto 0);
    signal conv34_1469 : std_logic_vector(7 downto 0);
    signal conv35x_xi_1248 : std_logic_vector(31 downto 0);
    signal conv39x_xi_1252 : std_logic_vector(31 downto 0);
    signal conv40_1479 : std_logic_vector(7 downto 0);
    signal conv46_1489 : std_logic_vector(7 downto 0);
    signal conv6_1419 : std_logic_vector(7 downto 0);
    signal conv89x_xi_1400 : std_logic_vector(7 downto 0);
    signal conv_1396 : std_logic_vector(63 downto 0);
    signal iNsTr_2_1220 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1278_delayed_1_0_1295 : std_logic_vector(31 downto 0);
    signal iNsTr_2_at_entry_1197 : std_logic_vector(31 downto 0);
    signal inc67x_xcolx_x1x_xi_1330 : std_logic_vector(15 downto 0);
    signal inc67x_xi_1322 : std_logic_vector(15 downto 0);
    signal inc76x_xi_1347 : std_logic_vector(15 downto 0);
    signal inc76x_xrow18x_x1x_xi_1355 : std_logic_vector(15 downto 0);
    signal inc76x_xrow18x_x1x_xix_xlcssa_1386 : std_logic_vector(15 downto 0);
    signal incx_xi_1312 : std_logic_vector(15 downto 0);
    signal mul40x_xi_1258 : std_logic_vector(31 downto 0);
    signal row18x_x1x_xi_1225 : std_logic_vector(15 downto 0);
    signal row18x_x1x_xi_1329_delayed_2_0_1350 : std_logic_vector(15 downto 0);
    signal row18x_x1x_xi_at_entry_1202 : std_logic_vector(15 downto 0);
    signal shlx_xi_1269 : std_logic_vector(31 downto 0);
    signal shr13_1435 : std_logic_vector(63 downto 0);
    signal shr19_1445 : std_logic_vector(63 downto 0);
    signal shr25_1455 : std_logic_vector(63 downto 0);
    signal shr31_1465 : std_logic_vector(63 downto 0);
    signal shr37_1475 : std_logic_vector(63 downto 0);
    signal shr43_1485 : std_logic_vector(63 downto 0);
    signal shr_1425 : std_logic_vector(63 downto 0);
    signal sub_1415 : std_logic_vector(63 downto 0);
    signal type_cast_1223_wire : std_logic_vector(31 downto 0);
    signal type_cast_1228_wire : std_logic_vector(15 downto 0);
    signal type_cast_1233_wire : std_logic_vector(15 downto 0);
    signal type_cast_1238_wire : std_logic_vector(15 downto 0);
    signal type_cast_1256_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1267_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1278_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1284_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1290_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1302_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1304_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1310_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1316_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1334_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1341_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1359_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1366_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1372_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1389_wire : std_logic_vector(15 downto 0);
    signal type_cast_1394_wire : std_logic_vector(63 downto 0);
    signal type_cast_1408_wire : std_logic_vector(63 downto 0);
    signal type_cast_1423_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1433_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1443_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1453_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1463_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1473_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1483_wire_constant : std_logic_vector(63 downto 0);
    signal whilex_xbodyx_xi_maxPool3Dx_xexit_taken_1377 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    chlx_x0x_xi_at_entry_1212 <= "0000000000000000";
    colx_x1x_xi_at_entry_1207 <= "0000000000000000";
    iNsTr_2_at_entry_1197 <= "00000000000000000000000000000000";
    row18x_x1x_xi_at_entry_1202 <= "0000000000000000";
    type_cast_1256_wire_constant <= "00000000000000000000000001110000";
    type_cast_1267_wire_constant <= "00000000000000000000000000000101";
    type_cast_1278_wire_constant <= "00000000000000000000000000010000";
    type_cast_1284_wire_constant <= "00000000000000000000011100000000";
    type_cast_1290_wire_constant <= "00000000000000000000011100010000";
    type_cast_1302_wire_constant <= "00000001";
    type_cast_1304_wire_constant <= "00000000";
    type_cast_1310_wire_constant <= "0000000000000001";
    type_cast_1316_wire_constant <= "0000000000010000";
    type_cast_1334_wire_constant <= "0000000000000000";
    type_cast_1341_wire_constant <= "0000000000111000";
    type_cast_1359_wire_constant <= "0000000000000000";
    type_cast_1366_wire_constant <= "00000000000000000000000000000001";
    type_cast_1372_wire_constant <= "0000000000111000";
    type_cast_1423_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1433_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1443_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1453_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1463_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1473_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1483_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    phi_stmt_1220: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1223_wire & iNsTr_2_at_entry_1197;
      req <= phi_stmt_1220_req_0 & phi_stmt_1220_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1220",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1220_ack_0,
          idata => idata,
          odata => iNsTr_2_1220,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1220
    phi_stmt_1225: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1228_wire & row18x_x1x_xi_at_entry_1202;
      req <= phi_stmt_1225_req_0 & phi_stmt_1225_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1225",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1225_ack_0,
          idata => idata,
          odata => row18x_x1x_xi_1225,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1225
    phi_stmt_1230: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1233_wire & colx_x1x_xi_at_entry_1207;
      req <= phi_stmt_1230_req_0 & phi_stmt_1230_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1230",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1230_ack_0,
          idata => idata,
          odata => colx_x1x_xi_1230,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1230
    phi_stmt_1235: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1238_wire & chlx_x0x_xi_at_entry_1212;
      req <= phi_stmt_1235_req_0 & phi_stmt_1235_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1235",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1235_ack_0,
          idata => idata,
          odata => chlx_x0x_xi_1235,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1235
    phi_stmt_1386: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1389_wire;
      req(0) <= phi_stmt_1386_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1386",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1386_ack_0,
          idata => idata,
          odata => inc76x_xrow18x_x1x_xix_xlcssa_1386,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1386
    -- flow-through select operator MUX_1336_inst
    chlx_x1x_xi_1337 <= type_cast_1334_wire_constant when (cmpx_xi_1318(0) /=  '0') else incx_xi_1312;
    -- flow-through select operator MUX_1361_inst
    colx_x2x_xi_1362 <= type_cast_1359_wire_constant when (cmp72x_xi_1343(0) /=  '0') else inc67x_xcolx_x1x_xi_1330;
    W_colx_x1x_xi_1307_delayed_1_0_1323_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_colx_x1x_xi_1307_delayed_1_0_1323_inst_req_0;
      W_colx_x1x_xi_1307_delayed_1_0_1323_inst_ack_0<= wack(0);
      rreq(0) <= W_colx_x1x_xi_1307_delayed_1_0_1323_inst_req_1;
      W_colx_x1x_xi_1307_delayed_1_0_1323_inst_ack_1<= rack(0);
      W_colx_x1x_xi_1307_delayed_1_0_1323_inst : InterlockBuffer generic map ( -- 
        name => "W_colx_x1x_xi_1307_delayed_1_0_1323_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => colx_x1x_xi_1230,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => colx_x1x_xi_1307_delayed_1_0_1325,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_iNsTr_2_1278_delayed_1_0_1293_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_iNsTr_2_1278_delayed_1_0_1293_inst_req_0;
      W_iNsTr_2_1278_delayed_1_0_1293_inst_ack_0<= wack(0);
      rreq(0) <= W_iNsTr_2_1278_delayed_1_0_1293_inst_req_1;
      W_iNsTr_2_1278_delayed_1_0_1293_inst_ack_1<= rack(0);
      W_iNsTr_2_1278_delayed_1_0_1293_inst : InterlockBuffer generic map ( -- 
        name => "W_iNsTr_2_1278_delayed_1_0_1293_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_2_1220,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_2_1278_delayed_1_0_1295,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_row18x_x1x_xi_1329_delayed_2_0_1348_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_row18x_x1x_xi_1329_delayed_2_0_1348_inst_req_0;
      W_row18x_x1x_xi_1329_delayed_2_0_1348_inst_ack_0<= wack(0);
      rreq(0) <= W_row18x_x1x_xi_1329_delayed_2_0_1348_inst_req_1;
      W_row18x_x1x_xi_1329_delayed_2_0_1348_inst_ack_1<= rack(0);
      W_row18x_x1x_xi_1329_delayed_2_0_1348_inst : InterlockBuffer generic map ( -- 
        name => "W_row18x_x1x_xi_1329_delayed_2_0_1348_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => row18x_x1x_xi_1225,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => row18x_x1x_xi_1329_delayed_2_0_1350,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_whilex_xbodyx_xi_maxPool3Dx_xexit_taken_1375_inst
    process(cmp84x_xi_1374) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := cmp84x_xi_1374(0 downto 0);
      whilex_xbodyx_xi_maxPool3Dx_xexit_taken_1377 <= tmp_var; -- 
    end process;
    type_cast_1223_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1223_inst_req_0;
      type_cast_1223_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1223_inst_req_1;
      type_cast_1223_inst_ack_1<= rack(0);
      type_cast_1223_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1223_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add79x_xi_1368,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1223_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1228_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1228_inst_req_0;
      type_cast_1228_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1228_inst_req_1;
      type_cast_1228_inst_ack_1<= rack(0);
      type_cast_1228_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1228_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc76x_xrow18x_x1x_xi_1355,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1228_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1233_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1233_inst_req_0;
      type_cast_1233_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1233_inst_req_1;
      type_cast_1233_inst_ack_1<= rack(0);
      type_cast_1233_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1233_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => colx_x2x_xi_1362,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1233_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1238_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1238_inst_req_0;
      type_cast_1238_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1238_inst_req_1;
      type_cast_1238_inst_ack_1<= rack(0);
      type_cast_1238_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1238_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => chlx_x1x_xi_1337,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1238_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1243_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1243_inst_req_0;
      type_cast_1243_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1243_inst_req_1;
      type_cast_1243_inst_ack_1<= rack(0);
      type_cast_1243_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1243_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => chlx_x0x_xi_1235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv31x_xi_1244,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1247_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1247_inst_req_0;
      type_cast_1247_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1247_inst_req_1;
      type_cast_1247_inst_ack_1<= rack(0);
      type_cast_1247_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1247_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => colx_x1x_xi_1230,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35x_xi_1248,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1251_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1251_inst_req_0;
      type_cast_1251_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1251_inst_req_1;
      type_cast_1251_inst_ack_1<= rack(0);
      type_cast_1251_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1251_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => row18x_x1x_xi_1225,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39x_xi_1252,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1321_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1321_inst_req_0;
      type_cast_1321_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1321_inst_req_1;
      type_cast_1321_inst_ack_1<= rack(0);
      type_cast_1321_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1321_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmpx_xi_1318,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc67x_xi_1322,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1346_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1346_inst_req_0;
      type_cast_1346_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1346_inst_req_1;
      type_cast_1346_inst_ack_1<= rack(0);
      type_cast_1346_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1346_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp72x_xi_1343,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc76x_xi_1347,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1389_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1389_inst_req_0;
      type_cast_1389_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1389_inst_req_1;
      type_cast_1389_inst_ack_1<= rack(0);
      type_cast_1389_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1389_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc76x_xrow18x_x1x_xi_1355,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1389_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1395_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1395_inst_req_0;
      type_cast_1395_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1395_inst_req_1;
      type_cast_1395_inst_ack_1<= rack(0);
      type_cast_1395_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1395_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1394_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1396,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1399_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1399_inst_req_0;
      type_cast_1399_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1399_inst_req_1;
      type_cast_1399_inst_ack_1<= rack(0);
      type_cast_1399_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1399_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc76x_xrow18x_x1x_xix_xlcssa_1386,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv89x_xi_1400,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1409_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1409_inst_req_0;
      type_cast_1409_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1409_inst_req_1;
      type_cast_1409_inst_ack_1<= rack(0);
      type_cast_1409_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1409_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1408_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2_1410,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1418_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1418_inst_req_0;
      type_cast_1418_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1418_inst_req_1;
      type_cast_1418_inst_ack_1<= rack(0);
      type_cast_1418_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1418_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_1415,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv6_1419,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1428_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1428_inst_req_0;
      type_cast_1428_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1428_inst_req_1;
      type_cast_1428_inst_ack_1<= rack(0);
      type_cast_1428_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1428_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_1425,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10_1429,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1438_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1438_inst_req_0;
      type_cast_1438_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1438_inst_req_1;
      type_cast_1438_inst_ack_1<= rack(0);
      type_cast_1438_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1438_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr13_1435,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv16_1439,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1448_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1448_inst_req_0;
      type_cast_1448_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1448_inst_req_1;
      type_cast_1448_inst_ack_1<= rack(0);
      type_cast_1448_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1448_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr19_1445,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_1449,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1458_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1458_inst_req_0;
      type_cast_1458_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1458_inst_req_1;
      type_cast_1458_inst_ack_1<= rack(0);
      type_cast_1458_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1458_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr25_1455,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv28_1459,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1468_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1468_inst_req_0;
      type_cast_1468_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1468_inst_req_1;
      type_cast_1468_inst_ack_1<= rack(0);
      type_cast_1468_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1468_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr31_1465,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv34_1469,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1478_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1478_inst_req_0;
      type_cast_1478_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1478_inst_req_1;
      type_cast_1478_inst_ack_1<= rack(0);
      type_cast_1478_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1478_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr37_1475,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv40_1479,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1488_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1488_inst_req_0;
      type_cast_1488_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1488_inst_req_1;
      type_cast_1488_inst_ack_1<= rack(0);
      type_cast_1488_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1488_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr43_1485,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv46_1489,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1218_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1380_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1218_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1218_branch_req_0,
          ack0 => do_while_stmt_1218_branch_ack_0,
          ack1 => do_while_stmt_1218_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1381_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= whilex_xbodyx_xi_maxPool3Dx_xexit_taken_1377;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1381_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1381_branch_req_0,
          ack0 => if_stmt_1381_branch_ack_0,
          ack1 => if_stmt_1381_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1311_inst
    process(chlx_x0x_xi_1235) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(chlx_x0x_xi_1235, type_cast_1310_wire_constant, tmp_var);
      incx_xi_1312 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1329_inst
    process(inc67x_xi_1322, colx_x1x_xi_1307_delayed_1_0_1325) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc67x_xi_1322, colx_x1x_xi_1307_delayed_1_0_1325, tmp_var);
      inc67x_xcolx_x1x_xi_1330 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1354_inst
    process(inc76x_xi_1347, row18x_x1x_xi_1329_delayed_2_0_1350) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc76x_xi_1347, row18x_x1x_xi_1329_delayed_2_0_1350, tmp_var);
      inc76x_xrow18x_x1x_xi_1355 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1262_inst
    process(conv35x_xi_1248, mul40x_xi_1258) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv35x_xi_1248, mul40x_xi_1258, tmp_var);
      add41x_xi_1263 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1273_inst
    process(shlx_xi_1269, conv31x_xi_1244) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shlx_xi_1269, conv31x_xi_1244, tmp_var);
      add43x_xi_1274 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1279_inst
    process(add43x_xi_1274) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add43x_xi_1274, type_cast_1278_wire_constant, tmp_var);
      add50x_xi_1280 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1285_inst
    process(add43x_xi_1274) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add43x_xi_1274, type_cast_1284_wire_constant, tmp_var);
      add54x_xi_1286 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1291_inst
    process(add43x_xi_1274) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add43x_xi_1274, type_cast_1290_wire_constant, tmp_var);
      add57x_xi_1292 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1367_inst
    process(iNsTr_2_1220) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_2_1220, type_cast_1366_wire_constant, tmp_var);
      add79x_xi_1368 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1317_inst
    process(incx_xi_1312) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(incx_xi_1312, type_cast_1316_wire_constant, tmp_var);
      cmpx_xi_1318 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1342_inst
    process(inc67x_xcolx_x1x_xi_1330) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc67x_xcolx_x1x_xi_1330, type_cast_1341_wire_constant, tmp_var);
      cmp72x_xi_1343 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1373_inst
    process(inc76x_xrow18x_x1x_xi_1355) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc76x_xrow18x_x1x_xi_1355, type_cast_1372_wire_constant, tmp_var);
      cmp84x_xi_1374 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1424_inst
    process(sub_1415) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1415, type_cast_1423_wire_constant, tmp_var);
      shr_1425 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1434_inst
    process(sub_1415) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1415, type_cast_1433_wire_constant, tmp_var);
      shr13_1435 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1444_inst
    process(sub_1415) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1415, type_cast_1443_wire_constant, tmp_var);
      shr19_1445 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1454_inst
    process(sub_1415) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1415, type_cast_1453_wire_constant, tmp_var);
      shr25_1455 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1464_inst
    process(sub_1415) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1415, type_cast_1463_wire_constant, tmp_var);
      shr31_1465 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1474_inst
    process(sub_1415) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1415, type_cast_1473_wire_constant, tmp_var);
      shr37_1475 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1484_inst
    process(sub_1415) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1415, type_cast_1483_wire_constant, tmp_var);
      shr43_1485 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1257_inst
    process(conv39x_xi_1252) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv39x_xi_1252, type_cast_1256_wire_constant, tmp_var);
      mul40x_xi_1258 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1380_inst
    process(cmp84x_xi_1374) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp84x_xi_1374, tmp_var);
      NOT_u1_u1_1380_wire <= tmp_var; -- 
    end process;
    -- binary operator SHL_u32_u32_1268_inst
    process(add41x_xi_1263) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add41x_xi_1263, type_cast_1267_wire_constant, tmp_var);
      shlx_xi_1269 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1414_inst
    process(conv2_1410, conv_1396) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv2_1410, conv_1396, tmp_var);
      sub_1415 <= tmp_var; --
    end process;
    -- unary operator type_cast_1394_inst
    process(call_1194) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call_1194, tmp_var);
      type_cast_1394_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1408_inst
    process(call1_1405) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call1_1405, tmp_var);
      type_cast_1408_wire <= tmp_var; -- 
    end process;
    -- shared outport operator group (0) : WPIPE_system_output_pipe_1490_inst WPIPE_system_output_pipe_1493_inst WPIPE_system_output_pipe_1511_inst WPIPE_system_output_pipe_1508_inst WPIPE_system_output_pipe_1401_inst WPIPE_system_output_pipe_1505_inst WPIPE_system_output_pipe_1502_inst WPIPE_system_output_pipe_1499_inst WPIPE_system_output_pipe_1496_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal sample_req, sample_ack : BooleanArray( 8 downto 0);
      signal update_req, update_ack : BooleanArray( 8 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 8 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 8 downto 0);
      signal guard_vector : std_logic_vector( 8 downto 0);
      constant inBUFs : IntegerArray(8 downto 0) := (8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(8 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false);
      constant guardBuffering: IntegerArray(8 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2);
      -- 
    begin -- 
      sample_req_unguarded(8) <= WPIPE_system_output_pipe_1490_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_system_output_pipe_1493_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_system_output_pipe_1511_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_system_output_pipe_1508_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_system_output_pipe_1401_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_system_output_pipe_1505_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_system_output_pipe_1502_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_system_output_pipe_1499_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_system_output_pipe_1496_inst_req_0;
      WPIPE_system_output_pipe_1490_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_system_output_pipe_1493_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_system_output_pipe_1511_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_system_output_pipe_1508_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_system_output_pipe_1401_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_system_output_pipe_1505_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_system_output_pipe_1502_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_system_output_pipe_1499_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_system_output_pipe_1496_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(8) <= WPIPE_system_output_pipe_1490_inst_req_1;
      update_req_unguarded(7) <= WPIPE_system_output_pipe_1493_inst_req_1;
      update_req_unguarded(6) <= WPIPE_system_output_pipe_1511_inst_req_1;
      update_req_unguarded(5) <= WPIPE_system_output_pipe_1508_inst_req_1;
      update_req_unguarded(4) <= WPIPE_system_output_pipe_1401_inst_req_1;
      update_req_unguarded(3) <= WPIPE_system_output_pipe_1505_inst_req_1;
      update_req_unguarded(2) <= WPIPE_system_output_pipe_1502_inst_req_1;
      update_req_unguarded(1) <= WPIPE_system_output_pipe_1499_inst_req_1;
      update_req_unguarded(0) <= WPIPE_system_output_pipe_1496_inst_req_1;
      WPIPE_system_output_pipe_1490_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_system_output_pipe_1493_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_system_output_pipe_1511_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_system_output_pipe_1508_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_system_output_pipe_1401_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_system_output_pipe_1505_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_system_output_pipe_1502_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_system_output_pipe_1499_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_system_output_pipe_1496_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      data_in <= conv46_1489 & conv40_1479 & conv6_1419 & conv10_1429 & conv89x_xi_1400 & conv16_1439 & conv22_1449 & conv28_1459 & conv34_1469;
      system_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "system_output_pipe_write_0_gI", nreqs => 9, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      system_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "system_output_pipe", data_width => 8, num_reqs => 9, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => system_output_pipe_pipe_write_req(0),
          oack => system_output_pipe_pipe_write_ack(0),
          odata => system_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1192_call 
    fill_input_call_group_0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1192_call_req_0;
      call_stmt_1192_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1192_call_req_1;
      call_stmt_1192_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      fill_input_call_group_0_gI: SplitGuardInterface generic map(name => "fill_input_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => fill_input_call_reqs(0),
          ackR => fill_input_call_acks(0),
          tagR => fill_input_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => fill_input_return_acks(0), -- cross-over
          ackL => fill_input_return_reqs(0), -- cross-over
          tagL => fill_input_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1405_call call_stmt_1194_call 
    timer_call_group_1: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1405_call_req_0;
      reqL_unguarded(0) <= call_stmt_1194_call_req_0;
      call_stmt_1405_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1194_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1405_call_req_1;
      reqR_unguarded(0) <= call_stmt_1194_call_req_1;
      call_stmt_1405_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1194_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_1_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_1_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_1_gI: SplitGuardInterface generic map(name => "timer_call_group_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call1_1405 <= data_out(127 downto 64);
      call_1194 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1306_call 
    maxPool4_call_group_2: Block -- 
      signal data_in: std_logic_vector(175 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 15);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1306_call_req_0;
      call_stmt_1306_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1306_call_req_1;
      call_stmt_1306_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      maxPool4_call_group_2_gI: SplitGuardInterface generic map(name => "maxPool4_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= iNsTr_2_1278_delayed_1_0_1295 & add43x_xi_1274 & add50x_xi_1280 & add54x_xi_1286 & add57x_xi_1292 & type_cast_1302_wire_constant & type_cast_1304_wire_constant;
      callx_xi_1306 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 176,
        owidth => 176,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => maxPool4_call_reqs(0),
          ackR => maxPool4_call_acks(0),
          dataR => maxPool4_call_data(175 downto 0),
          tagR => maxPool4_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => maxPool4_return_acks(0), -- cross-over
          ackL => maxPool4_return_reqs(0), -- cross-over
          dataL => maxPool4_return_data(7 downto 0),
          tagL => maxPool4_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_1514_call 
    sendOutput_call_group_3: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1514_call_req_0;
      call_stmt_1514_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1514_call_req_1;
      call_stmt_1514_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendOutput_call_group_3_gI: SplitGuardInterface generic map(name => "sendOutput_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => sendOutput_call_reqs(0),
          ackR => sendOutput_call_acks(0),
          tagR => sendOutput_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendOutput_return_acks(0), -- cross-over
          ackL => sendOutput_return_reqs(0), -- cross-over
          tagL => sendOutput_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- 
  end Block; -- data_path
  -- 
end systemTOP_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    T : out  std_logic_vector(63 downto 0);
    timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
    timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal T_buffer :  std_logic_vector(63 downto 0);
  signal T_update_enable: Boolean;
  signal timer_CP_2011_start: Boolean;
  signal timer_CP_2011_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_req_1182_inst_req_0 : boolean;
  signal WPIPE_timer_req_1182_inst_ack_0 : boolean;
  signal WPIPE_timer_req_1182_inst_req_1 : boolean;
  signal WPIPE_timer_req_1182_inst_ack_1 : boolean;
  signal RPIPE_timer_resp_1187_inst_req_0 : boolean;
  signal RPIPE_timer_resp_1187_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_1187_inst_req_1 : boolean;
  signal RPIPE_timer_resp_1187_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_2011_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= T_buffer;
  T <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_2011_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_2011_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_2011_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_2011: Block -- control-path 
    signal timer_CP_2011_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    timer_CP_2011_elements(0) <= timer_CP_2011_start;
    timer_CP_2011_symbol <= timer_CP_2011_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_1185_to_assign_stmt_1188/$entry
      -- CP-element group 0: 	 assign_stmt_1185_to_assign_stmt_1188/WPIPE_timer_req_1182_sample_start_
      -- CP-element group 0: 	 assign_stmt_1185_to_assign_stmt_1188/WPIPE_timer_req_1182_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1185_to_assign_stmt_1188/WPIPE_timer_req_1182_Sample/req
      -- CP-element group 0: 	 assign_stmt_1185_to_assign_stmt_1188/RPIPE_timer_resp_1187_sample_start_
      -- CP-element group 0: 	 assign_stmt_1185_to_assign_stmt_1188/RPIPE_timer_resp_1187_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1185_to_assign_stmt_1188/RPIPE_timer_resp_1187_Sample/rr
      -- 
    rr_2038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_2011_elements(0), ack => RPIPE_timer_resp_1187_inst_req_0); -- 
    req_2024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_2011_elements(0), ack => WPIPE_timer_req_1182_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_1185_to_assign_stmt_1188/WPIPE_timer_req_1182_sample_completed_
      -- CP-element group 1: 	 assign_stmt_1185_to_assign_stmt_1188/WPIPE_timer_req_1182_update_start_
      -- CP-element group 1: 	 assign_stmt_1185_to_assign_stmt_1188/WPIPE_timer_req_1182_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1185_to_assign_stmt_1188/WPIPE_timer_req_1182_Sample/ack
      -- CP-element group 1: 	 assign_stmt_1185_to_assign_stmt_1188/WPIPE_timer_req_1182_Update/$entry
      -- CP-element group 1: 	 assign_stmt_1185_to_assign_stmt_1188/WPIPE_timer_req_1182_Update/req
      -- 
    ack_2025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_1182_inst_ack_0, ack => timer_CP_2011_elements(1)); -- 
    req_2029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_2011_elements(1), ack => WPIPE_timer_req_1182_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_1185_to_assign_stmt_1188/WPIPE_timer_req_1182_update_completed_
      -- CP-element group 2: 	 assign_stmt_1185_to_assign_stmt_1188/WPIPE_timer_req_1182_Update/$exit
      -- CP-element group 2: 	 assign_stmt_1185_to_assign_stmt_1188/WPIPE_timer_req_1182_Update/ack
      -- 
    ack_2030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_1182_inst_ack_1, ack => timer_CP_2011_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_1185_to_assign_stmt_1188/RPIPE_timer_resp_1187_sample_completed_
      -- CP-element group 3: 	 assign_stmt_1185_to_assign_stmt_1188/RPIPE_timer_resp_1187_update_start_
      -- CP-element group 3: 	 assign_stmt_1185_to_assign_stmt_1188/RPIPE_timer_resp_1187_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_1185_to_assign_stmt_1188/RPIPE_timer_resp_1187_Sample/ra
      -- CP-element group 3: 	 assign_stmt_1185_to_assign_stmt_1188/RPIPE_timer_resp_1187_Update/$entry
      -- CP-element group 3: 	 assign_stmt_1185_to_assign_stmt_1188/RPIPE_timer_resp_1187_Update/cr
      -- 
    ra_2039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_1187_inst_ack_0, ack => timer_CP_2011_elements(3)); -- 
    cr_2043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_2011_elements(3), ack => RPIPE_timer_resp_1187_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_1185_to_assign_stmt_1188/RPIPE_timer_resp_1187_update_completed_
      -- CP-element group 4: 	 assign_stmt_1185_to_assign_stmt_1188/RPIPE_timer_resp_1187_Update/$exit
      -- CP-element group 4: 	 assign_stmt_1185_to_assign_stmt_1188/RPIPE_timer_resp_1187_Update/ca
      -- 
    ca_2044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_1187_inst_ack_1, ack => timer_CP_2011_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_1185_to_assign_stmt_1188/$exit
      -- 
    timer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "timer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timer_CP_2011_elements(2) & timer_CP_2011_elements(4);
      gj_timer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timer_CP_2011_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal type_cast_1184_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_1184_wire_constant <= "1";
    -- shared inport operator group (0) : RPIPE_timer_resp_1187_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_resp_1187_inst_req_0;
      RPIPE_timer_resp_1187_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_resp_1187_inst_req_1;
      RPIPE_timer_resp_1187_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      T_buffer <= data_out(63 downto 0);
      timer_resp_read_0_gI: SplitGuardInterface generic map(name => "timer_resp_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_resp_read_0: InputPortRevised -- 
        generic map ( name => "timer_resp_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_resp_pipe_read_req(0),
          oack => timer_resp_pipe_read_ack(0),
          odata => timer_resp_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_req_1182_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_req_1182_inst_req_0;
      WPIPE_timer_req_1182_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_req_1182_inst_req_1;
      WPIPE_timer_req_1182_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1184_wire_constant;
      timer_req_write_0_gI: SplitGuardInterface generic map(name => "timer_req_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_req_write_0: OutputPortRevised -- 
        generic map ( name => "timer_req", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_req_pipe_write_req(0),
          oack => timer_req_pipe_write_ack(0),
          odata => timer_req_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_2809_start: Boolean;
  signal timerDaemon_CP_2809_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal nCOUNTER_1536_1527_buf_ack_0 : boolean;
  signal phi_stmt_1523_req_1 : boolean;
  signal nCOUNTER_1536_1527_buf_req_1 : boolean;
  signal nCOUNTER_1536_1527_buf_ack_1 : boolean;
  signal nCOUNTER_1536_1527_buf_req_0 : boolean;
  signal phi_stmt_1523_ack_0 : boolean;
  signal do_while_stmt_1521_branch_req_0 : boolean;
  signal phi_stmt_1523_req_0 : boolean;
  signal RPIPE_timer_req_1530_inst_req_0 : boolean;
  signal RPIPE_timer_req_1530_inst_ack_0 : boolean;
  signal RPIPE_timer_req_1530_inst_req_1 : boolean;
  signal RPIPE_timer_req_1530_inst_ack_1 : boolean;
  signal WPIPE_timer_resp_1538_inst_req_0 : boolean;
  signal WPIPE_timer_resp_1538_inst_ack_0 : boolean;
  signal WPIPE_timer_resp_1538_inst_req_1 : boolean;
  signal WPIPE_timer_resp_1538_inst_ack_1 : boolean;
  signal do_while_stmt_1521_branch_ack_0 : boolean;
  signal do_while_stmt_1521_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_2809_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_2809_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_2809_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_2809_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_2809: Block -- control-path 
    signal timerDaemon_CP_2809_elements: BooleanArray(44 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_2809_elements(0) <= timerDaemon_CP_2809_start;
    timerDaemon_CP_2809_symbol <= timerDaemon_CP_2809_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1520/$entry
      -- CP-element group 0: 	 branch_block_stmt_1520/do_while_stmt_1521__entry__
      -- CP-element group 0: 	 branch_block_stmt_1520/branch_block_stmt_1520__entry__
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	44 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1520/$exit
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1520/branch_block_stmt_1520__exit__
      -- CP-element group 1: 	 branch_block_stmt_1520/do_while_stmt_1521__exit__
      -- 
    timerDaemon_CP_2809_elements(1) <= timerDaemon_CP_2809_elements(44);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1520/do_while_stmt_1521/$entry
      -- CP-element group 2: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521__entry__
      -- 
    timerDaemon_CP_2809_elements(2) <= timerDaemon_CP_2809_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	44 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521__exit__
      -- 
    -- Element group timerDaemon_CP_2809_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1520/do_while_stmt_1521/loop_back
      -- 
    -- Element group timerDaemon_CP_2809_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	42 
    -- CP-element group 5: 	43 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1520/do_while_stmt_1521/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1520/do_while_stmt_1521/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1520/do_while_stmt_1521/loop_taken/$entry
      -- 
    timerDaemon_CP_2809_elements(5) <= timerDaemon_CP_2809_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	41 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1520/do_while_stmt_1521/loop_body_done
      -- 
    timerDaemon_CP_2809_elements(6) <= timerDaemon_CP_2809_elements(41);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_2809_elements(7) <= timerDaemon_CP_2809_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_2809_elements(8) <= timerDaemon_CP_2809_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	40 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/phi_stmt_1528_sample_start_
      -- 
    -- Element group timerDaemon_CP_2809_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	40 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/condition_evaluated
      -- 
    condition_evaluated_2833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2809_elements(10), ack => do_while_stmt_1521_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2809_elements(14) & timerDaemon_CP_2809_elements(40);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2809_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/phi_stmt_1523_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_2809_elements(9) & timerDaemon_CP_2809_elements(15) & timerDaemon_CP_2809_elements(14);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2809_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	41 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/phi_stmt_1523_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/phi_stmt_1528_sample_completed_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2809_elements(17) & timerDaemon_CP_2809_elements(35);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2809_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	32 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/phi_stmt_1523_update_start__ps
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2809_elements(16) & timerDaemon_CP_2809_elements(32);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2809_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/aggregated_phi_update_ack
      -- 
    timerDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2809_elements(18) & timerDaemon_CP_2809_elements(36);
      gj_timerDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2809_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/phi_stmt_1523_sample_start_
      -- 
    timerDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2809_elements(9) & timerDaemon_CP_2809_elements(12);
      gj_timerDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2809_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	38 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/phi_stmt_1523_update_start_
      -- 
    timerDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2809_elements(9) & timerDaemon_CP_2809_elements(38);
      gj_timerDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2809_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/phi_stmt_1523_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_2809_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	37 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/phi_stmt_1523_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/phi_stmt_1523_update_completed_
      -- 
    -- Element group timerDaemon_CP_2809_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/phi_stmt_1523_loopback_trigger
      -- 
    timerDaemon_CP_2809_elements(19) <= timerDaemon_CP_2809_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/phi_stmt_1523_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/phi_stmt_1523_loopback_sample_req_ps
      -- 
    phi_stmt_1523_loopback_sample_req_2848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1523_loopback_sample_req_2848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2809_elements(20), ack => phi_stmt_1523_req_1); -- 
    -- Element group timerDaemon_CP_2809_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/phi_stmt_1523_entry_trigger
      -- 
    timerDaemon_CP_2809_elements(21) <= timerDaemon_CP_2809_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/phi_stmt_1523_entry_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/phi_stmt_1523_entry_sample_req
      -- 
    phi_stmt_1523_entry_sample_req_2851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1523_entry_sample_req_2851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2809_elements(22), ack => phi_stmt_1523_req_0); -- 
    -- Element group timerDaemon_CP_2809_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/phi_stmt_1523_phi_mux_ack_ps
      -- CP-element group 23: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/phi_stmt_1523_phi_mux_ack
      -- 
    phi_stmt_1523_phi_mux_ack_2854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1523_ack_0, ack => timerDaemon_CP_2809_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/type_cast_1526_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/type_cast_1526_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/type_cast_1526_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/type_cast_1526_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_2809_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/type_cast_1526_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/type_cast_1526_update_start_
      -- 
    -- Element group timerDaemon_CP_2809_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/type_cast_1526_update_completed__ps
      -- 
    timerDaemon_CP_2809_elements(26) <= timerDaemon_CP_2809_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/type_cast_1526_update_completed_
      -- 
    -- Element group timerDaemon_CP_2809_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => timerDaemon_CP_2809_elements(25), ack => timerDaemon_CP_2809_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/R_nCOUNTER_1527_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/R_nCOUNTER_1527_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/R_nCOUNTER_1527_Sample/req
      -- CP-element group 28: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/R_nCOUNTER_1527_Sample/$entry
      -- 
    req_2875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2809_elements(28), ack => nCOUNTER_1536_1527_buf_req_0); -- 
    -- Element group timerDaemon_CP_2809_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/R_nCOUNTER_1527_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/R_nCOUNTER_1527_Update/req
      -- CP-element group 29: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/R_nCOUNTER_1527_update_start_
      -- CP-element group 29: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/R_nCOUNTER_1527_Update/$entry
      -- 
    req_2880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2809_elements(29), ack => nCOUNTER_1536_1527_buf_req_1); -- 
    -- Element group timerDaemon_CP_2809_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/R_nCOUNTER_1527_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/R_nCOUNTER_1527_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/R_nCOUNTER_1527_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/R_nCOUNTER_1527_Sample/$exit
      -- 
    ack_2876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_1536_1527_buf_ack_0, ack => timerDaemon_CP_2809_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/R_nCOUNTER_1527_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/R_nCOUNTER_1527_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/R_nCOUNTER_1527_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/R_nCOUNTER_1527_update_completed_
      -- 
    ack_2881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_1536_1527_buf_ack_1, ack => timerDaemon_CP_2809_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	38 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/phi_stmt_1528_update_start_
      -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2809_elements(9) & timerDaemon_CP_2809_elements(38);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2809_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/RPIPE_timer_req_1530_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/RPIPE_timer_req_1530_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/RPIPE_timer_req_1530_Sample/rr
      -- 
    rr_2894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2809_elements(33), ack => RPIPE_timer_req_1530_inst_req_0); -- 
    timerDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2809_elements(11) & timerDaemon_CP_2809_elements(36);
      gj_timerDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2809_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/RPIPE_timer_req_1530_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/RPIPE_timer_req_1530_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/RPIPE_timer_req_1530_Update/cr
      -- 
    cr_2899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2809_elements(34), ack => RPIPE_timer_req_1530_inst_req_1); -- 
    timerDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2809_elements(13) & timerDaemon_CP_2809_elements(35);
      gj_timerDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2809_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/RPIPE_timer_req_1530_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/RPIPE_timer_req_1530_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/RPIPE_timer_req_1530_Sample/ra
      -- 
    ra_2895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_1530_inst_ack_0, ack => timerDaemon_CP_2809_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	37 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/phi_stmt_1528_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/RPIPE_timer_req_1530_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/RPIPE_timer_req_1530_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/RPIPE_timer_req_1530_Update/ca
      -- 
    ca_2900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_1530_inst_ack_1, ack => timerDaemon_CP_2809_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	18 
    -- CP-element group 37: 	36 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/WPIPE_timer_resp_1538_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/WPIPE_timer_resp_1538_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/WPIPE_timer_resp_1538_Sample/req
      -- 
    req_2908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2809_elements(37), ack => WPIPE_timer_resp_1538_inst_req_0); -- 
    timerDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_2809_elements(18) & timerDaemon_CP_2809_elements(36) & timerDaemon_CP_2809_elements(39);
      gj_timerDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2809_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	16 
    -- CP-element group 38: 	32 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/WPIPE_timer_resp_1538_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/WPIPE_timer_resp_1538_update_start_
      -- CP-element group 38: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/WPIPE_timer_resp_1538_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/WPIPE_timer_resp_1538_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/WPIPE_timer_resp_1538_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/WPIPE_timer_resp_1538_Update/req
      -- 
    ack_2909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_1538_inst_ack_0, ack => timerDaemon_CP_2809_elements(38)); -- 
    req_2913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2809_elements(38), ack => WPIPE_timer_resp_1538_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/WPIPE_timer_resp_1538_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/WPIPE_timer_resp_1538_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/WPIPE_timer_resp_1538_Update/ack
      -- 
    ack_2914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_1538_inst_ack_1, ack => timerDaemon_CP_2809_elements(39)); -- 
    -- CP-element group 40:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	10 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_2809_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => timerDaemon_CP_2809_elements(9), ack => timerDaemon_CP_2809_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	12 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	6 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1520/do_while_stmt_1521/do_while_stmt_1521_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2809_elements(12) & timerDaemon_CP_2809_elements(39);
      gj_timerDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2809_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	5 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1520/do_while_stmt_1521/loop_exit/$exit
      -- CP-element group 42: 	 branch_block_stmt_1520/do_while_stmt_1521/loop_exit/ack
      -- 
    ack_2919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1521_branch_ack_0, ack => timerDaemon_CP_2809_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	5 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1520/do_while_stmt_1521/loop_taken/$exit
      -- CP-element group 43: 	 branch_block_stmt_1520/do_while_stmt_1521/loop_taken/ack
      -- 
    ack_2923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1521_branch_ack_1, ack => timerDaemon_CP_2809_elements(43)); -- 
    -- CP-element group 44:  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	3 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	1 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_1520/do_while_stmt_1521/$exit
      -- 
    timerDaemon_CP_2809_elements(44) <= timerDaemon_CP_2809_elements(3);
    timerDaemon_do_while_stmt_1521_terminator_2924: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_1521_terminator_2924", max_iterations_in_flight =>7) 
      port map(loop_body_exit => timerDaemon_CP_2809_elements(6),loop_continue => timerDaemon_CP_2809_elements(43),loop_terminate => timerDaemon_CP_2809_elements(42),loop_back => timerDaemon_CP_2809_elements(4),loop_exit => timerDaemon_CP_2809_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1523_phi_seq_2882_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_2809_elements(21);
      timerDaemon_CP_2809_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_2809_elements(24);
      timerDaemon_CP_2809_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_2809_elements(26);
      timerDaemon_CP_2809_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_2809_elements(19);
      timerDaemon_CP_2809_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_2809_elements(30);
      timerDaemon_CP_2809_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_2809_elements(31);
      timerDaemon_CP_2809_elements(20) <= phi_mux_reqs(1);
      phi_stmt_1523_phi_seq_2882 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1523_phi_seq_2882") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_2809_elements(11), 
          phi_sample_ack => timerDaemon_CP_2809_elements(17), 
          phi_update_req => timerDaemon_CP_2809_elements(13), 
          phi_update_ack => timerDaemon_CP_2809_elements(18), 
          phi_mux_ack => timerDaemon_CP_2809_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2834_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_2809_elements(7);
        preds(1)  <= timerDaemon_CP_2809_elements(8);
        entry_tmerge_2834 : transition_merge -- 
          generic map(name => " entry_tmerge_2834")
          port map (preds => preds, symbol_out => timerDaemon_CP_2809_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal COUNTER_1523 : std_logic_vector(63 downto 0);
    signal RPIPE_timer_req_1530_wire : std_logic_vector(0 downto 0);
    signal konst_1534_wire_constant : std_logic_vector(63 downto 0);
    signal konst_1542_wire_constant : std_logic_vector(0 downto 0);
    signal nCOUNTER_1536 : std_logic_vector(63 downto 0);
    signal nCOUNTER_1536_1527_buffered : std_logic_vector(63 downto 0);
    signal req_1528 : std_logic_vector(0 downto 0);
    signal type_cast_1526_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_1534_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_1542_wire_constant <= "1";
    type_cast_1526_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_1523: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1526_wire_constant & nCOUNTER_1536_1527_buffered;
      req <= phi_stmt_1523_req_0 & phi_stmt_1523_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1523",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1523_ack_0,
          idata => idata,
          odata => COUNTER_1523,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1523
    nCOUNTER_1536_1527_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nCOUNTER_1536_1527_buf_req_0;
      nCOUNTER_1536_1527_buf_ack_0<= wack(0);
      rreq(0) <= nCOUNTER_1536_1527_buf_req_1;
      nCOUNTER_1536_1527_buf_ack_1<= rack(0);
      nCOUNTER_1536_1527_buf : InterlockBuffer generic map ( -- 
        name => "nCOUNTER_1536_1527_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nCOUNTER_1536,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nCOUNTER_1536_1527_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_1528
    process(RPIPE_timer_req_1530_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := RPIPE_timer_req_1530_wire(0 downto 0);
      req_1528 <= tmp_var; -- 
    end process;
    do_while_stmt_1521_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1542_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1521_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1521_branch_req_0,
          ack0 => do_while_stmt_1521_branch_ack_0,
          ack1 => do_while_stmt_1521_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_1535_inst
    process(COUNTER_1523) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(COUNTER_1523, konst_1534_wire_constant, tmp_var);
      nCOUNTER_1536 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_timer_req_1530_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_req_1530_inst_req_0;
      RPIPE_timer_req_1530_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_req_1530_inst_req_1;
      RPIPE_timer_req_1530_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_timer_req_1530_wire <= data_out(0 downto 0);
      timer_req_read_0_gI: SplitGuardInterface generic map(name => "timer_req_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_req_read_0: InputPortRevised -- 
        generic map ( name => "timer_req_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_req_pipe_read_req(0),
          oack => timer_req_pipe_read_ack(0),
          odata => timer_req_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_resp_1538_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_resp_1538_inst_req_0;
      WPIPE_timer_resp_1538_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_resp_1538_inst_req_1;
      WPIPE_timer_resp_1538_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= req_1528(0);
      data_in <= COUNTER_1523;
      timer_resp_write_0_gI: SplitGuardInterface generic map(name => "timer_resp_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_resp_write_0: OutputPortRevised -- 
        generic map ( name => "timer_resp", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_resp_pipe_write_req(0),
          oack => timer_resp_pipe_write_ack(0),
          odata => timer_resp_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity writeModule1 is -- 
  generic (tag_length : integer); 
  port ( -- 
    address : in  std_logic_vector(31 downto 0);
    data : in  std_logic_vector(63 downto 0);
    memoryModule_call_reqs : out  std_logic_vector(0 downto 0);
    memoryModule_call_acks : in   std_logic_vector(0 downto 0);
    memoryModule_call_data : out  std_logic_vector(96 downto 0);
    memoryModule_call_tag  :  out  std_logic_vector(0 downto 0);
    memoryModule_return_reqs : out  std_logic_vector(0 downto 0);
    memoryModule_return_acks : in   std_logic_vector(0 downto 0);
    memoryModule_return_data : in   std_logic_vector(63 downto 0);
    memoryModule_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writeModule1;
architecture writeModule1_arch of writeModule1 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 96)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal address_buffer :  std_logic_vector(31 downto 0);
  signal address_update_enable: Boolean;
  signal data_buffer :  std_logic_vector(63 downto 0);
  signal data_update_enable: Boolean;
  -- output port buffer signals
  signal writeModule1_CP_102_start: Boolean;
  signal writeModule1_CP_102_symbol: Boolean;
  -- volatile/operator module components. 
  component memoryModule is -- 
    generic (tag_length : integer); 
    port ( -- 
      r_wbar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(31 downto 0);
      data_in : in  std_logic_vector(63 downto 0);
      data_out : out  std_logic_vector(63 downto 0);
      MAIN_MEM_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MAIN_MEM_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MAIN_MEM_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      MAIN_MEM_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      MAIN_MEM_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      MAIN_MEM_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_70_call_req_0 : boolean;
  signal call_stmt_70_call_ack_0 : boolean;
  signal call_stmt_70_call_req_1 : boolean;
  signal call_stmt_70_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writeModule1_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 96) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= address;
  address_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(95 downto 32) <= data;
  data_buffer <= in_buffer_data_out(95 downto 32);
  in_buffer_data_in(tag_length + 95 downto 96) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 95 downto 96);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writeModule1_CP_102_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writeModule1_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeModule1_CP_102_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writeModule1_CP_102_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeModule1_CP_102_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writeModule1_CP_102: Block -- control-path 
    signal writeModule1_CP_102_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    writeModule1_CP_102_elements(0) <= writeModule1_CP_102_start;
    writeModule1_CP_102_symbol <= writeModule1_CP_102_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_70/$entry
      -- CP-element group 0: 	 call_stmt_70/call_stmt_70_sample_start_
      -- CP-element group 0: 	 call_stmt_70/call_stmt_70_update_start_
      -- CP-element group 0: 	 call_stmt_70/call_stmt_70_Sample/$entry
      -- CP-element group 0: 	 call_stmt_70/call_stmt_70_Sample/crr
      -- CP-element group 0: 	 call_stmt_70/call_stmt_70_Update/$entry
      -- CP-element group 0: 	 call_stmt_70/call_stmt_70_Update/ccr
      -- 
    crr_115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_102_elements(0), ack => call_stmt_70_call_req_0); -- 
    ccr_120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_102_elements(0), ack => call_stmt_70_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_70/call_stmt_70_sample_completed_
      -- CP-element group 1: 	 call_stmt_70/call_stmt_70_Sample/$exit
      -- CP-element group 1: 	 call_stmt_70/call_stmt_70_Sample/cra
      -- 
    cra_116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_70_call_ack_0, ack => writeModule1_CP_102_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_70/$exit
      -- CP-element group 2: 	 call_stmt_70/call_stmt_70_update_completed_
      -- CP-element group 2: 	 call_stmt_70/call_stmt_70_Update/$exit
      -- CP-element group 2: 	 call_stmt_70/call_stmt_70_Update/cca
      -- 
    cca_121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_70_call_ack_1, ack => writeModule1_CP_102_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_67_wire : std_logic_vector(31 downto 0);
    signal konst_64_wire_constant : std_logic_vector(0 downto 0);
    signal konst_65_wire_constant : std_logic_vector(31 downto 0);
    signal out1_70 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_64_wire_constant <= "0";
    konst_65_wire_constant <= "00000000000000000000000000000000";
    -- binary operator ADD_u32_u32_67_inst
    process(address_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address_buffer, konst_65_wire_constant, tmp_var);
      ADD_u32_u32_67_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_70_call 
    memoryModule_call_group_0: Block -- 
      signal data_in: std_logic_vector(96 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_70_call_req_0;
      call_stmt_70_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_70_call_req_1;
      call_stmt_70_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      memoryModule_call_group_0_gI: SplitGuardInterface generic map(name => "memoryModule_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_64_wire_constant & ADD_u32_u32_67_wire & data_buffer;
      out1_70 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 97,
        owidth => 97,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => memoryModule_call_reqs(0),
          ackR => memoryModule_call_acks(0),
          dataR => memoryModule_call_data(96 downto 0),
          tagR => memoryModule_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => memoryModule_return_acks(0), -- cross-over
          ackL => memoryModule_return_reqs(0), -- cross-over
          dataL => memoryModule_return_data(63 downto 0),
          tagL => memoryModule_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writeModule1_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity writeModule_maxPool is -- 
  generic (tag_length : integer); 
  port ( -- 
    index : in  std_logic_vector(7 downto 0);
    address : in  std_logic_vector(31 downto 0);
    data : in  std_logic_vector(63 downto 0);
    done : out  std_logic_vector(0 downto 0);
    memoryModule_call_reqs : out  std_logic_vector(0 downto 0);
    memoryModule_call_acks : in   std_logic_vector(0 downto 0);
    memoryModule_call_data : out  std_logic_vector(96 downto 0);
    memoryModule_call_tag  :  out  std_logic_vector(0 downto 0);
    memoryModule_return_reqs : out  std_logic_vector(0 downto 0);
    memoryModule_return_acks : in   std_logic_vector(0 downto 0);
    memoryModule_return_data : in   std_logic_vector(63 downto 0);
    memoryModule_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writeModule_maxPool;
architecture writeModule_maxPool_arch of writeModule_maxPool is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 104)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal index_buffer :  std_logic_vector(7 downto 0);
  signal index_update_enable: Boolean;
  signal address_buffer :  std_logic_vector(31 downto 0);
  signal address_update_enable: Boolean;
  signal data_buffer :  std_logic_vector(63 downto 0);
  signal data_update_enable: Boolean;
  -- output port buffer signals
  signal done_buffer :  std_logic_vector(0 downto 0);
  signal done_update_enable: Boolean;
  signal writeModule_maxPool_CP_517_start: Boolean;
  signal writeModule_maxPool_CP_517_symbol: Boolean;
  -- volatile/operator module components. 
  component memoryModule is -- 
    generic (tag_length : integer); 
    port ( -- 
      r_wbar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(31 downto 0);
      data_in : in  std_logic_vector(63 downto 0);
      data_out : out  std_logic_vector(63 downto 0);
      MAIN_MEM_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MAIN_MEM_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MAIN_MEM_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      MAIN_MEM_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      MAIN_MEM_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      MAIN_MEM_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal BITSEL_u8_u1_278_inst_ack_1 : boolean;
  signal BITSEL_u8_u1_278_inst_req_1 : boolean;
  signal BITSEL_u8_u1_278_inst_ack_0 : boolean;
  signal BITSEL_u8_u1_278_inst_req_0 : boolean;
  signal call_stmt_274_call_ack_1 : boolean;
  signal call_stmt_274_call_req_1 : boolean;
  signal call_stmt_274_call_ack_0 : boolean;
  signal call_stmt_274_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writeModule_maxPool_input_buffer", -- 
      buffer_size => 2,
      bypass_flag => false,
      data_width => tag_length + 104) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= index;
  index_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(39 downto 8) <= address;
  address_buffer <= in_buffer_data_out(39 downto 8);
  in_buffer_data_in(103 downto 40) <= data;
  data_buffer <= in_buffer_data_out(103 downto 40);
  in_buffer_data_in(tag_length + 103 downto 104) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 103 downto 104);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 4) := (0 => 8,1 => 8,2 => 8,3 => 1,4 => 8);
    constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 8);
    constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 5); -- 
  begin -- 
    preds <= index_update_enable & address_update_enable & data_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writeModule_maxPool_CP_517_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writeModule_maxPool_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= done_buffer;
  done <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 8);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeModule_maxPool_CP_517_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  done_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 23) := "done_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_done_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => done_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 8,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writeModule_maxPool_CP_517_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeModule_maxPool_CP_517_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writeModule_maxPool_CP_517: Block -- control-path 
    signal writeModule_maxPool_CP_517_elements: BooleanArray(19 downto 0);
    -- 
  begin -- 
    writeModule_maxPool_CP_517_elements(0) <= writeModule_maxPool_CP_517_start;
    writeModule_maxPool_CP_517_symbol <= writeModule_maxPool_CP_517_elements(19);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	10 
    -- CP-element group 1: 	6 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 call_stmt_274_to_assign_stmt_279/$entry
      -- 
    writeModule_maxPool_CP_517_elements(1) <= writeModule_maxPool_CP_517_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	12 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	15 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 call_stmt_274_to_assign_stmt_279/index_update_enable
      -- CP-element group 2: 	 call_stmt_274_to_assign_stmt_279/index_update_enable_out
      -- 
    writeModule_maxPool_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "writeModule_maxPool_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeModule_maxPool_CP_517_elements(12);
      gj_writeModule_maxPool_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule_maxPool_CP_517_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	8 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	16 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 call_stmt_274_to_assign_stmt_279/address_update_enable
      -- CP-element group 3: 	 call_stmt_274_to_assign_stmt_279/address_update_enable_out
      -- 
    writeModule_maxPool_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "writeModule_maxPool_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeModule_maxPool_CP_517_elements(8);
      gj_writeModule_maxPool_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule_maxPool_CP_517_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	8 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	17 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 call_stmt_274_to_assign_stmt_279/data_update_enable_out
      -- CP-element group 4: 	 call_stmt_274_to_assign_stmt_279/data_update_enable
      -- 
    writeModule_maxPool_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "writeModule_maxPool_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeModule_maxPool_CP_517_elements(8);
      gj_writeModule_maxPool_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule_maxPool_CP_517_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	18 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	11 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 call_stmt_274_to_assign_stmt_279/done_update_enable_in
      -- CP-element group 5: 	 call_stmt_274_to_assign_stmt_279/done_update_enable
      -- 
    writeModule_maxPool_CP_517_elements(5) <= writeModule_maxPool_CP_517_elements(18);
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	1 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	8 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 call_stmt_274_to_assign_stmt_279/call_stmt_274_Sample/$entry
      -- CP-element group 6: 	 call_stmt_274_to_assign_stmt_279/call_stmt_274_sample_start_
      -- CP-element group 6: 	 call_stmt_274_to_assign_stmt_279/call_stmt_274_Sample/crr
      -- 
    crr_538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule_maxPool_CP_517_elements(6), ack => call_stmt_274_call_req_0); -- 
    writeModule_maxPool_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "writeModule_maxPool_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule_maxPool_CP_517_elements(1) & writeModule_maxPool_CP_517_elements(8);
      gj_writeModule_maxPool_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule_maxPool_CP_517_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: marked-predecessors 
    -- CP-element group 7: 	9 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	9 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_274_to_assign_stmt_279/call_stmt_274_update_start_
      -- CP-element group 7: 	 call_stmt_274_to_assign_stmt_279/call_stmt_274_Update/ccr
      -- CP-element group 7: 	 call_stmt_274_to_assign_stmt_279/call_stmt_274_Update/$entry
      -- 
    ccr_543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule_maxPool_CP_517_elements(7), ack => call_stmt_274_call_req_1); -- 
    writeModule_maxPool_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "writeModule_maxPool_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeModule_maxPool_CP_517_elements(9);
      gj_writeModule_maxPool_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule_maxPool_CP_517_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: 	3 
    -- CP-element group 8: 	4 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_274_to_assign_stmt_279/call_stmt_274_sample_completed_
      -- CP-element group 8: 	 call_stmt_274_to_assign_stmt_279/call_stmt_274_Sample/cra
      -- CP-element group 8: 	 call_stmt_274_to_assign_stmt_279/call_stmt_274_Sample/$exit
      -- 
    cra_539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_274_call_ack_0, ack => writeModule_maxPool_CP_517_elements(8)); -- 
    -- CP-element group 9:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	7 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	14 
    -- CP-element group 9: marked-successors 
    -- CP-element group 9: 	7 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 call_stmt_274_to_assign_stmt_279/call_stmt_274_update_completed_
      -- CP-element group 9: 	 call_stmt_274_to_assign_stmt_279/call_stmt_274_Update/cca
      -- CP-element group 9: 	 call_stmt_274_to_assign_stmt_279/call_stmt_274_Update/$exit
      -- 
    cca_544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_274_call_ack_1, ack => writeModule_maxPool_CP_517_elements(9)); -- 
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	1 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_274_to_assign_stmt_279/BITSEL_u8_u1_278_Sample/rr
      -- CP-element group 10: 	 call_stmt_274_to_assign_stmt_279/BITSEL_u8_u1_278_Sample/$entry
      -- CP-element group 10: 	 call_stmt_274_to_assign_stmt_279/BITSEL_u8_u1_278_sample_start_
      -- 
    rr_552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule_maxPool_CP_517_elements(10), ack => BITSEL_u8_u1_278_inst_req_0); -- 
    writeModule_maxPool_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "writeModule_maxPool_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule_maxPool_CP_517_elements(1) & writeModule_maxPool_CP_517_elements(12);
      gj_writeModule_maxPool_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule_maxPool_CP_517_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	5 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	13 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_274_to_assign_stmt_279/BITSEL_u8_u1_278_Update/cr
      -- CP-element group 11: 	 call_stmt_274_to_assign_stmt_279/BITSEL_u8_u1_278_Update/$entry
      -- CP-element group 11: 	 call_stmt_274_to_assign_stmt_279/BITSEL_u8_u1_278_update_start_
      -- 
    cr_557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule_maxPool_CP_517_elements(11), ack => BITSEL_u8_u1_278_inst_req_1); -- 
    writeModule_maxPool_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "writeModule_maxPool_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule_maxPool_CP_517_elements(5) & writeModule_maxPool_CP_517_elements(13);
      gj_writeModule_maxPool_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule_maxPool_CP_517_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: 	2 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_274_to_assign_stmt_279/BITSEL_u8_u1_278_Sample/ra
      -- CP-element group 12: 	 call_stmt_274_to_assign_stmt_279/BITSEL_u8_u1_278_Sample/$exit
      -- CP-element group 12: 	 call_stmt_274_to_assign_stmt_279/BITSEL_u8_u1_278_sample_completed_
      -- 
    ra_553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => BITSEL_u8_u1_278_inst_ack_0, ack => writeModule_maxPool_CP_517_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	11 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_274_to_assign_stmt_279/BITSEL_u8_u1_278_update_completed_
      -- CP-element group 13: 	 call_stmt_274_to_assign_stmt_279/BITSEL_u8_u1_278_Update/ca
      -- CP-element group 13: 	 call_stmt_274_to_assign_stmt_279/BITSEL_u8_u1_278_Update/$exit
      -- 
    ca_558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => BITSEL_u8_u1_278_inst_ack_1, ack => writeModule_maxPool_CP_517_elements(13)); -- 
    -- CP-element group 14:  join  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	9 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	19 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 call_stmt_274_to_assign_stmt_279/$exit
      -- 
    writeModule_maxPool_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 8);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "writeModule_maxPool_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule_maxPool_CP_517_elements(9) & writeModule_maxPool_CP_517_elements(13);
      gj_writeModule_maxPool_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule_maxPool_CP_517_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 index_update_enable
      -- 
    writeModule_maxPool_CP_517_elements(15) <= writeModule_maxPool_CP_517_elements(2);
    -- CP-element group 16:  place  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	3 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 address_update_enable
      -- 
    writeModule_maxPool_CP_517_elements(16) <= writeModule_maxPool_CP_517_elements(3);
    -- CP-element group 17:  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	4 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 data_update_enable
      -- 
    writeModule_maxPool_CP_517_elements(17) <= writeModule_maxPool_CP_517_elements(4);
    -- CP-element group 18:  place  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	5 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 done_update_enable
      -- 
    -- CP-element group 19:  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	14 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 $exit
      -- 
    writeModule_maxPool_CP_517_elements(19) <= writeModule_maxPool_CP_517_elements(14);
    --  hookup: inputs to control-path 
    writeModule_maxPool_CP_517_elements(18) <= done_update_enable;
    -- hookup: output from control-path 
    data_update_enable <= writeModule_maxPool_CP_517_elements(17);
    address_update_enable <= writeModule_maxPool_CP_517_elements(16);
    index_update_enable <= writeModule_maxPool_CP_517_elements(15);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_271_wire : std_logic_vector(31 downto 0);
    signal konst_268_wire_constant : std_logic_vector(0 downto 0);
    signal konst_269_wire_constant : std_logic_vector(31 downto 0);
    signal konst_277_wire_constant : std_logic_vector(7 downto 0);
    signal out1_274 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_268_wire_constant <= "0";
    konst_269_wire_constant <= "00000000000000000000000000000000";
    konst_277_wire_constant <= "00000000";
    -- binary operator ADD_u32_u32_271_inst
    process(address_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address_buffer, konst_269_wire_constant, tmp_var);
      ADD_u32_u32_271_wire <= tmp_var; --
    end process;
    -- shared split operator group (1) : BITSEL_u8_u1_278_inst 
    ApBitsel_group_1: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= index_buffer;
      done_buffer <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= BITSEL_u8_u1_278_inst_req_0;
      BITSEL_u8_u1_278_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= BITSEL_u8_u1_278_inst_req_1;
      BITSEL_u8_u1_278_inst_ack_1 <= ackR_unguarded(0);
      ApBitsel_group_1_gI: SplitGuardInterface generic map(name => "ApBitsel_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApBitsel",
          name => "ApBitsel_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared call operator group (0) : call_stmt_274_call 
    memoryModule_call_group_0: Block -- 
      signal data_in: std_logic_vector(96 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_274_call_req_0;
      call_stmt_274_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_274_call_req_1;
      call_stmt_274_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      memoryModule_call_group_0_gI: SplitGuardInterface generic map(name => "memoryModule_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_268_wire_constant & ADD_u32_u32_271_wire & data_buffer;
      out1_274 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 97,
        owidth => 97,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => memoryModule_call_reqs(0),
          ackR => memoryModule_call_acks(0),
          dataR => memoryModule_call_data(96 downto 0),
          tagR => memoryModule_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => memoryModule_return_acks(0), -- cross-over
          ackL => memoryModule_return_reqs(0), -- cross-over
          dataL => memoryModule_return_data(63 downto 0),
          tagL => memoryModule_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writeModule_maxPool_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    MAIN_MEM_REQUEST_pipe_read_data: out std_logic_vector(109 downto 0);
    MAIN_MEM_REQUEST_pipe_read_req : in std_logic_vector(0 downto 0);
    MAIN_MEM_REQUEST_pipe_read_ack : out std_logic_vector(0 downto 0);
    MAIN_MEM_RESPONSE_pipe_write_data: in std_logic_vector(64 downto 0);
    MAIN_MEM_RESPONSE_pipe_write_req : in std_logic_vector(0 downto 0);
    MAIN_MEM_RESPONSE_pipe_write_ack : out std_logic_vector(0 downto 0);
    system_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    system_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    system_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    system_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    system_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    system_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- declarations related to module fill_input
  component fill_input is -- 
    generic (tag_length : integer); 
    port ( -- 
      system_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      system_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      system_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      writeModule1_call_reqs : out  std_logic_vector(0 downto 0);
      writeModule1_call_acks : in   std_logic_vector(0 downto 0);
      writeModule1_call_data : out  std_logic_vector(95 downto 0);
      writeModule1_call_tag  :  out  std_logic_vector(0 downto 0);
      writeModule1_return_reqs : out  std_logic_vector(0 downto 0);
      writeModule1_return_acks : in   std_logic_vector(0 downto 0);
      writeModule1_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module fill_input
  signal fill_input_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal fill_input_tag_out   : std_logic_vector(1 downto 0);
  signal fill_input_start_req : std_logic;
  signal fill_input_start_ack : std_logic;
  signal fill_input_fin_req   : std_logic;
  signal fill_input_fin_ack : std_logic;
  -- caller side aggregated signals for module fill_input
  signal fill_input_call_reqs: std_logic_vector(0 downto 0);
  signal fill_input_call_acks: std_logic_vector(0 downto 0);
  signal fill_input_return_reqs: std_logic_vector(0 downto 0);
  signal fill_input_return_acks: std_logic_vector(0 downto 0);
  signal fill_input_call_tag: std_logic_vector(0 downto 0);
  signal fill_input_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module maxPool4
  component maxPool4 is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(31 downto 0);
      addr1 : in  std_logic_vector(31 downto 0);
      addr2 : in  std_logic_vector(31 downto 0);
      addr3 : in  std_logic_vector(31 downto 0);
      addr4 : in  std_logic_vector(31 downto 0);
      index1 : in  std_logic_vector(7 downto 0);
      index2 : in  std_logic_vector(7 downto 0);
      output : out  std_logic_vector(7 downto 0);
      readModule_maxPool_call_reqs : out  std_logic_vector(0 downto 0);
      readModule_maxPool_call_acks : in   std_logic_vector(0 downto 0);
      readModule_maxPool_call_data : out  std_logic_vector(39 downto 0);
      readModule_maxPool_call_tag  :  out  std_logic_vector(2 downto 0);
      readModule_maxPool_return_reqs : out  std_logic_vector(0 downto 0);
      readModule_maxPool_return_acks : in   std_logic_vector(0 downto 0);
      readModule_maxPool_return_data : in   std_logic_vector(63 downto 0);
      readModule_maxPool_return_tag :  in   std_logic_vector(2 downto 0);
      writeModule_maxPool_call_reqs : out  std_logic_vector(0 downto 0);
      writeModule_maxPool_call_acks : in   std_logic_vector(0 downto 0);
      writeModule_maxPool_call_data : out  std_logic_vector(103 downto 0);
      writeModule_maxPool_call_tag  :  out  std_logic_vector(0 downto 0);
      writeModule_maxPool_return_reqs : out  std_logic_vector(0 downto 0);
      writeModule_maxPool_return_acks : in   std_logic_vector(0 downto 0);
      writeModule_maxPool_return_data : in   std_logic_vector(0 downto 0);
      writeModule_maxPool_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module maxPool4
  signal maxPool4_addr :  std_logic_vector(31 downto 0);
  signal maxPool4_addr1 :  std_logic_vector(31 downto 0);
  signal maxPool4_addr2 :  std_logic_vector(31 downto 0);
  signal maxPool4_addr3 :  std_logic_vector(31 downto 0);
  signal maxPool4_addr4 :  std_logic_vector(31 downto 0);
  signal maxPool4_index1 :  std_logic_vector(7 downto 0);
  signal maxPool4_index2 :  std_logic_vector(7 downto 0);
  signal maxPool4_output :  std_logic_vector(7 downto 0);
  signal maxPool4_in_args    : std_logic_vector(175 downto 0);
  signal maxPool4_out_args   : std_logic_vector(7 downto 0);
  signal maxPool4_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal maxPool4_tag_out   : std_logic_vector(1 downto 0);
  signal maxPool4_start_req : std_logic;
  signal maxPool4_start_ack : std_logic;
  signal maxPool4_fin_req   : std_logic;
  signal maxPool4_fin_ack : std_logic;
  -- caller side aggregated signals for module maxPool4
  signal maxPool4_call_reqs: std_logic_vector(0 downto 0);
  signal maxPool4_call_acks: std_logic_vector(0 downto 0);
  signal maxPool4_return_reqs: std_logic_vector(0 downto 0);
  signal maxPool4_return_acks: std_logic_vector(0 downto 0);
  signal maxPool4_call_data: std_logic_vector(175 downto 0);
  signal maxPool4_call_tag: std_logic_vector(0 downto 0);
  signal maxPool4_return_data: std_logic_vector(7 downto 0);
  signal maxPool4_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module memoryModule
  component memoryModule is -- 
    generic (tag_length : integer); 
    port ( -- 
      r_wbar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(31 downto 0);
      data_in : in  std_logic_vector(63 downto 0);
      data_out : out  std_logic_vector(63 downto 0);
      MAIN_MEM_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MAIN_MEM_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MAIN_MEM_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      MAIN_MEM_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      MAIN_MEM_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      MAIN_MEM_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module memoryModule
  signal memoryModule_r_wbar :  std_logic_vector(0 downto 0);
  signal memoryModule_addr :  std_logic_vector(31 downto 0);
  signal memoryModule_data_in :  std_logic_vector(63 downto 0);
  signal memoryModule_data_out :  std_logic_vector(63 downto 0);
  signal memoryModule_in_args    : std_logic_vector(96 downto 0);
  signal memoryModule_out_args   : std_logic_vector(63 downto 0);
  signal memoryModule_tag_in    : std_logic_vector(3 downto 0) := (others => '0');
  signal memoryModule_tag_out   : std_logic_vector(3 downto 0);
  signal memoryModule_start_req : std_logic;
  signal memoryModule_start_ack : std_logic;
  signal memoryModule_fin_req   : std_logic;
  signal memoryModule_fin_ack : std_logic;
  -- caller side aggregated signals for module memoryModule
  signal memoryModule_call_reqs: std_logic_vector(3 downto 0);
  signal memoryModule_call_acks: std_logic_vector(3 downto 0);
  signal memoryModule_return_reqs: std_logic_vector(3 downto 0);
  signal memoryModule_return_acks: std_logic_vector(3 downto 0);
  signal memoryModule_call_data: std_logic_vector(387 downto 0);
  signal memoryModule_call_tag: std_logic_vector(3 downto 0);
  signal memoryModule_return_data: std_logic_vector(255 downto 0);
  signal memoryModule_return_tag: std_logic_vector(3 downto 0);
  -- declarations related to module readModule1
  component readModule1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      address : in  std_logic_vector(31 downto 0);
      data : out  std_logic_vector(63 downto 0);
      memoryModule_call_reqs : out  std_logic_vector(0 downto 0);
      memoryModule_call_acks : in   std_logic_vector(0 downto 0);
      memoryModule_call_data : out  std_logic_vector(96 downto 0);
      memoryModule_call_tag  :  out  std_logic_vector(0 downto 0);
      memoryModule_return_reqs : out  std_logic_vector(0 downto 0);
      memoryModule_return_acks : in   std_logic_vector(0 downto 0);
      memoryModule_return_data : in   std_logic_vector(63 downto 0);
      memoryModule_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module readModule1
  signal readModule1_address :  std_logic_vector(31 downto 0);
  signal readModule1_data :  std_logic_vector(63 downto 0);
  signal readModule1_in_args    : std_logic_vector(31 downto 0);
  signal readModule1_out_args   : std_logic_vector(63 downto 0);
  signal readModule1_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal readModule1_tag_out   : std_logic_vector(1 downto 0);
  signal readModule1_start_req : std_logic;
  signal readModule1_start_ack : std_logic;
  signal readModule1_fin_req   : std_logic;
  signal readModule1_fin_ack : std_logic;
  -- caller side aggregated signals for module readModule1
  signal readModule1_call_reqs: std_logic_vector(0 downto 0);
  signal readModule1_call_acks: std_logic_vector(0 downto 0);
  signal readModule1_return_reqs: std_logic_vector(0 downto 0);
  signal readModule1_return_acks: std_logic_vector(0 downto 0);
  signal readModule1_call_data: std_logic_vector(31 downto 0);
  signal readModule1_call_tag: std_logic_vector(0 downto 0);
  signal readModule1_return_data: std_logic_vector(63 downto 0);
  signal readModule1_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module readModule_maxPool
  component readModule_maxPool is -- 
    generic (tag_length : integer); 
    port ( -- 
      index : in  std_logic_vector(7 downto 0);
      address : in  std_logic_vector(31 downto 0);
      data : out  std_logic_vector(63 downto 0);
      memoryModule_call_reqs : out  std_logic_vector(0 downto 0);
      memoryModule_call_acks : in   std_logic_vector(0 downto 0);
      memoryModule_call_data : out  std_logic_vector(96 downto 0);
      memoryModule_call_tag  :  out  std_logic_vector(0 downto 0);
      memoryModule_return_reqs : out  std_logic_vector(0 downto 0);
      memoryModule_return_acks : in   std_logic_vector(0 downto 0);
      memoryModule_return_data : in   std_logic_vector(63 downto 0);
      memoryModule_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module readModule_maxPool
  signal readModule_maxPool_index :  std_logic_vector(7 downto 0);
  signal readModule_maxPool_address :  std_logic_vector(31 downto 0);
  signal readModule_maxPool_data :  std_logic_vector(63 downto 0);
  signal readModule_maxPool_in_args    : std_logic_vector(39 downto 0);
  signal readModule_maxPool_out_args   : std_logic_vector(63 downto 0);
  signal readModule_maxPool_tag_in    : std_logic_vector(3 downto 0) := (others => '0');
  signal readModule_maxPool_tag_out   : std_logic_vector(3 downto 0);
  signal readModule_maxPool_start_req : std_logic;
  signal readModule_maxPool_start_ack : std_logic;
  signal readModule_maxPool_fin_req   : std_logic;
  signal readModule_maxPool_fin_ack : std_logic;
  -- caller side aggregated signals for module readModule_maxPool
  signal readModule_maxPool_call_reqs: std_logic_vector(0 downto 0);
  signal readModule_maxPool_call_acks: std_logic_vector(0 downto 0);
  signal readModule_maxPool_return_reqs: std_logic_vector(0 downto 0);
  signal readModule_maxPool_return_acks: std_logic_vector(0 downto 0);
  signal readModule_maxPool_call_data: std_logic_vector(39 downto 0);
  signal readModule_maxPool_call_tag: std_logic_vector(2 downto 0);
  signal readModule_maxPool_return_data: std_logic_vector(63 downto 0);
  signal readModule_maxPool_return_tag: std_logic_vector(2 downto 0);
  -- declarations related to module sendOutput
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      system_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      system_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      system_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      readModule1_call_reqs : out  std_logic_vector(0 downto 0);
      readModule1_call_acks : in   std_logic_vector(0 downto 0);
      readModule1_call_data : out  std_logic_vector(31 downto 0);
      readModule1_call_tag  :  out  std_logic_vector(0 downto 0);
      readModule1_return_reqs : out  std_logic_vector(0 downto 0);
      readModule1_return_acks : in   std_logic_vector(0 downto 0);
      readModule1_return_data : in   std_logic_vector(63 downto 0);
      readModule1_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendOutput
  signal sendOutput_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendOutput_tag_out   : std_logic_vector(1 downto 0);
  signal sendOutput_start_req : std_logic;
  signal sendOutput_start_ack : std_logic;
  signal sendOutput_fin_req   : std_logic;
  signal sendOutput_fin_ack : std_logic;
  -- caller side aggregated signals for module sendOutput
  signal sendOutput_call_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_call_acks: std_logic_vector(0 downto 0);
  signal sendOutput_return_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_return_acks: std_logic_vector(0 downto 0);
  signal sendOutput_call_tag: std_logic_vector(0 downto 0);
  signal sendOutput_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module systemTOP
  component systemTOP is -- 
    generic (tag_length : integer); 
    port ( -- 
      system_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      system_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      system_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      fill_input_call_reqs : out  std_logic_vector(0 downto 0);
      fill_input_call_acks : in   std_logic_vector(0 downto 0);
      fill_input_call_tag  :  out  std_logic_vector(0 downto 0);
      fill_input_return_reqs : out  std_logic_vector(0 downto 0);
      fill_input_return_acks : in   std_logic_vector(0 downto 0);
      fill_input_return_tag :  in   std_logic_vector(0 downto 0);
      maxPool4_call_reqs : out  std_logic_vector(0 downto 0);
      maxPool4_call_acks : in   std_logic_vector(0 downto 0);
      maxPool4_call_data : out  std_logic_vector(175 downto 0);
      maxPool4_call_tag  :  out  std_logic_vector(0 downto 0);
      maxPool4_return_reqs : out  std_logic_vector(0 downto 0);
      maxPool4_return_acks : in   std_logic_vector(0 downto 0);
      maxPool4_return_data : in   std_logic_vector(7 downto 0);
      maxPool4_return_tag :  in   std_logic_vector(0 downto 0);
      sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_call_acks : in   std_logic_vector(0 downto 0);
      sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
      sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_return_acks : in   std_logic_vector(0 downto 0);
      sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module systemTOP
  signal systemTOP_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal systemTOP_tag_out   : std_logic_vector(1 downto 0);
  signal systemTOP_start_req : std_logic;
  signal systemTOP_start_ack : std_logic;
  signal systemTOP_fin_req   : std_logic;
  signal systemTOP_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_T :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- declarations related to module writeModule1
  component writeModule1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      address : in  std_logic_vector(31 downto 0);
      data : in  std_logic_vector(63 downto 0);
      memoryModule_call_reqs : out  std_logic_vector(0 downto 0);
      memoryModule_call_acks : in   std_logic_vector(0 downto 0);
      memoryModule_call_data : out  std_logic_vector(96 downto 0);
      memoryModule_call_tag  :  out  std_logic_vector(0 downto 0);
      memoryModule_return_reqs : out  std_logic_vector(0 downto 0);
      memoryModule_return_acks : in   std_logic_vector(0 downto 0);
      memoryModule_return_data : in   std_logic_vector(63 downto 0);
      memoryModule_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writeModule1
  signal writeModule1_address :  std_logic_vector(31 downto 0);
  signal writeModule1_data :  std_logic_vector(63 downto 0);
  signal writeModule1_in_args    : std_logic_vector(95 downto 0);
  signal writeModule1_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writeModule1_tag_out   : std_logic_vector(1 downto 0);
  signal writeModule1_start_req : std_logic;
  signal writeModule1_start_ack : std_logic;
  signal writeModule1_fin_req   : std_logic;
  signal writeModule1_fin_ack : std_logic;
  -- caller side aggregated signals for module writeModule1
  signal writeModule1_call_reqs: std_logic_vector(0 downto 0);
  signal writeModule1_call_acks: std_logic_vector(0 downto 0);
  signal writeModule1_return_reqs: std_logic_vector(0 downto 0);
  signal writeModule1_return_acks: std_logic_vector(0 downto 0);
  signal writeModule1_call_data: std_logic_vector(95 downto 0);
  signal writeModule1_call_tag: std_logic_vector(0 downto 0);
  signal writeModule1_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module writeModule_maxPool
  component writeModule_maxPool is -- 
    generic (tag_length : integer); 
    port ( -- 
      index : in  std_logic_vector(7 downto 0);
      address : in  std_logic_vector(31 downto 0);
      data : in  std_logic_vector(63 downto 0);
      done : out  std_logic_vector(0 downto 0);
      memoryModule_call_reqs : out  std_logic_vector(0 downto 0);
      memoryModule_call_acks : in   std_logic_vector(0 downto 0);
      memoryModule_call_data : out  std_logic_vector(96 downto 0);
      memoryModule_call_tag  :  out  std_logic_vector(0 downto 0);
      memoryModule_return_reqs : out  std_logic_vector(0 downto 0);
      memoryModule_return_acks : in   std_logic_vector(0 downto 0);
      memoryModule_return_data : in   std_logic_vector(63 downto 0);
      memoryModule_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writeModule_maxPool
  signal writeModule_maxPool_index :  std_logic_vector(7 downto 0);
  signal writeModule_maxPool_address :  std_logic_vector(31 downto 0);
  signal writeModule_maxPool_data :  std_logic_vector(63 downto 0);
  signal writeModule_maxPool_done :  std_logic_vector(0 downto 0);
  signal writeModule_maxPool_in_args    : std_logic_vector(103 downto 0);
  signal writeModule_maxPool_out_args   : std_logic_vector(0 downto 0);
  signal writeModule_maxPool_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writeModule_maxPool_tag_out   : std_logic_vector(1 downto 0);
  signal writeModule_maxPool_start_req : std_logic;
  signal writeModule_maxPool_start_ack : std_logic;
  signal writeModule_maxPool_fin_req   : std_logic;
  signal writeModule_maxPool_fin_ack : std_logic;
  -- caller side aggregated signals for module writeModule_maxPool
  signal writeModule_maxPool_call_reqs: std_logic_vector(0 downto 0);
  signal writeModule_maxPool_call_acks: std_logic_vector(0 downto 0);
  signal writeModule_maxPool_return_reqs: std_logic_vector(0 downto 0);
  signal writeModule_maxPool_return_acks: std_logic_vector(0 downto 0);
  signal writeModule_maxPool_call_data: std_logic_vector(103 downto 0);
  signal writeModule_maxPool_call_tag: std_logic_vector(0 downto 0);
  signal writeModule_maxPool_return_data: std_logic_vector(0 downto 0);
  signal writeModule_maxPool_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe MAIN_MEM_REQUEST
  signal MAIN_MEM_REQUEST_pipe_write_data: std_logic_vector(109 downto 0);
  signal MAIN_MEM_REQUEST_pipe_write_req: std_logic_vector(0 downto 0);
  signal MAIN_MEM_REQUEST_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe MAIN_MEM_RESPONSE
  signal MAIN_MEM_RESPONSE_pipe_read_data: std_logic_vector(64 downto 0);
  signal MAIN_MEM_RESPONSE_pipe_read_req: std_logic_vector(0 downto 0);
  signal MAIN_MEM_RESPONSE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe system_input_pipe
  signal system_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal system_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal system_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe system_output_pipe
  signal system_output_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal system_output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal system_output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe timer_req
  signal timer_req_pipe_write_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_req
  signal timer_req_pipe_read_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_resp
  signal timer_resp_pipe_write_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_resp
  signal timer_resp_pipe_read_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module fill_input
  -- call arbiter for module fill_input
  fill_input_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => fill_input_call_reqs,
      call_acks => fill_input_call_acks,
      return_reqs => fill_input_return_reqs,
      return_acks => fill_input_return_acks,
      call_tag  => fill_input_call_tag,
      return_tag  => fill_input_return_tag,
      call_mtag => fill_input_tag_in,
      return_mtag => fill_input_tag_out,
      call_mreq => fill_input_start_req,
      call_mack => fill_input_start_ack,
      return_mreq => fill_input_fin_req,
      return_mack => fill_input_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  fill_input_instance:fill_input-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => fill_input_start_req,
      start_ack => fill_input_start_ack,
      fin_req => fill_input_fin_req,
      fin_ack => fill_input_fin_ack,
      clk => clk,
      reset => reset,
      system_input_pipe_pipe_read_req => system_input_pipe_pipe_read_req(0 downto 0),
      system_input_pipe_pipe_read_ack => system_input_pipe_pipe_read_ack(0 downto 0),
      system_input_pipe_pipe_read_data => system_input_pipe_pipe_read_data(7 downto 0),
      writeModule1_call_reqs => writeModule1_call_reqs(0 downto 0),
      writeModule1_call_acks => writeModule1_call_acks(0 downto 0),
      writeModule1_call_data => writeModule1_call_data(95 downto 0),
      writeModule1_call_tag => writeModule1_call_tag(0 downto 0),
      writeModule1_return_reqs => writeModule1_return_reqs(0 downto 0),
      writeModule1_return_acks => writeModule1_return_acks(0 downto 0),
      writeModule1_return_tag => writeModule1_return_tag(0 downto 0),
      tag_in => fill_input_tag_in,
      tag_out => fill_input_tag_out-- 
    ); -- 
  -- module maxPool4
  maxPool4_addr <= maxPool4_in_args(175 downto 144);
  maxPool4_addr1 <= maxPool4_in_args(143 downto 112);
  maxPool4_addr2 <= maxPool4_in_args(111 downto 80);
  maxPool4_addr3 <= maxPool4_in_args(79 downto 48);
  maxPool4_addr4 <= maxPool4_in_args(47 downto 16);
  maxPool4_index1 <= maxPool4_in_args(15 downto 8);
  maxPool4_index2 <= maxPool4_in_args(7 downto 0);
  maxPool4_out_args <= maxPool4_output ;
  -- call arbiter for module maxPool4
  maxPool4_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 176,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => maxPool4_call_reqs,
      call_acks => maxPool4_call_acks,
      return_reqs => maxPool4_return_reqs,
      return_acks => maxPool4_return_acks,
      call_data  => maxPool4_call_data,
      call_tag  => maxPool4_call_tag,
      return_tag  => maxPool4_return_tag,
      call_mtag => maxPool4_tag_in,
      return_mtag => maxPool4_tag_out,
      return_data =>maxPool4_return_data,
      call_mreq => maxPool4_start_req,
      call_mack => maxPool4_start_ack,
      return_mreq => maxPool4_fin_req,
      return_mack => maxPool4_fin_ack,
      call_mdata => maxPool4_in_args,
      return_mdata => maxPool4_out_args,
      clk => clk, 
      reset => reset --
    ); --
  maxPool4_instance:maxPool4-- 
    generic map(tag_length => 2)
    port map(-- 
      addr => maxPool4_addr,
      addr1 => maxPool4_addr1,
      addr2 => maxPool4_addr2,
      addr3 => maxPool4_addr3,
      addr4 => maxPool4_addr4,
      index1 => maxPool4_index1,
      index2 => maxPool4_index2,
      output => maxPool4_output,
      start_req => maxPool4_start_req,
      start_ack => maxPool4_start_ack,
      fin_req => maxPool4_fin_req,
      fin_ack => maxPool4_fin_ack,
      clk => clk,
      reset => reset,
      readModule_maxPool_call_reqs => readModule_maxPool_call_reqs(0 downto 0),
      readModule_maxPool_call_acks => readModule_maxPool_call_acks(0 downto 0),
      readModule_maxPool_call_data => readModule_maxPool_call_data(39 downto 0),
      readModule_maxPool_call_tag => readModule_maxPool_call_tag(2 downto 0),
      readModule_maxPool_return_reqs => readModule_maxPool_return_reqs(0 downto 0),
      readModule_maxPool_return_acks => readModule_maxPool_return_acks(0 downto 0),
      readModule_maxPool_return_data => readModule_maxPool_return_data(63 downto 0),
      readModule_maxPool_return_tag => readModule_maxPool_return_tag(2 downto 0),
      writeModule_maxPool_call_reqs => writeModule_maxPool_call_reqs(0 downto 0),
      writeModule_maxPool_call_acks => writeModule_maxPool_call_acks(0 downto 0),
      writeModule_maxPool_call_data => writeModule_maxPool_call_data(103 downto 0),
      writeModule_maxPool_call_tag => writeModule_maxPool_call_tag(0 downto 0),
      writeModule_maxPool_return_reqs => writeModule_maxPool_return_reqs(0 downto 0),
      writeModule_maxPool_return_acks => writeModule_maxPool_return_acks(0 downto 0),
      writeModule_maxPool_return_data => writeModule_maxPool_return_data(0 downto 0),
      writeModule_maxPool_return_tag => writeModule_maxPool_return_tag(0 downto 0),
      tag_in => maxPool4_tag_in,
      tag_out => maxPool4_tag_out-- 
    ); -- 
  -- module memoryModule
  memoryModule_r_wbar <= memoryModule_in_args(96 downto 96);
  memoryModule_addr <= memoryModule_in_args(95 downto 64);
  memoryModule_data_in <= memoryModule_in_args(63 downto 0);
  memoryModule_out_args <= memoryModule_data_out ;
  -- call arbiter for module memoryModule
  memoryModule_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 4,
      call_data_width => 97,
      return_data_width => 64,
      callee_tag_length => 3,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => memoryModule_call_reqs,
      call_acks => memoryModule_call_acks,
      return_reqs => memoryModule_return_reqs,
      return_acks => memoryModule_return_acks,
      call_data  => memoryModule_call_data,
      call_tag  => memoryModule_call_tag,
      return_tag  => memoryModule_return_tag,
      call_mtag => memoryModule_tag_in,
      return_mtag => memoryModule_tag_out,
      return_data =>memoryModule_return_data,
      call_mreq => memoryModule_start_req,
      call_mack => memoryModule_start_ack,
      return_mreq => memoryModule_fin_req,
      return_mack => memoryModule_fin_ack,
      call_mdata => memoryModule_in_args,
      return_mdata => memoryModule_out_args,
      clk => clk, 
      reset => reset --
    ); --
  memoryModule_instance:memoryModule-- 
    generic map(tag_length => 4)
    port map(-- 
      r_wbar => memoryModule_r_wbar,
      addr => memoryModule_addr,
      data_in => memoryModule_data_in,
      data_out => memoryModule_data_out,
      start_req => memoryModule_start_req,
      start_ack => memoryModule_start_ack,
      fin_req => memoryModule_fin_req,
      fin_ack => memoryModule_fin_ack,
      clk => clk,
      reset => reset,
      MAIN_MEM_RESPONSE_pipe_read_req => MAIN_MEM_RESPONSE_pipe_read_req(0 downto 0),
      MAIN_MEM_RESPONSE_pipe_read_ack => MAIN_MEM_RESPONSE_pipe_read_ack(0 downto 0),
      MAIN_MEM_RESPONSE_pipe_read_data => MAIN_MEM_RESPONSE_pipe_read_data(64 downto 0),
      MAIN_MEM_REQUEST_pipe_write_req => MAIN_MEM_REQUEST_pipe_write_req(0 downto 0),
      MAIN_MEM_REQUEST_pipe_write_ack => MAIN_MEM_REQUEST_pipe_write_ack(0 downto 0),
      MAIN_MEM_REQUEST_pipe_write_data => MAIN_MEM_REQUEST_pipe_write_data(109 downto 0),
      tag_in => memoryModule_tag_in,
      tag_out => memoryModule_tag_out-- 
    ); -- 
  -- module readModule1
  readModule1_address <= readModule1_in_args(31 downto 0);
  readModule1_out_args <= readModule1_data ;
  -- call arbiter for module readModule1
  readModule1_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 32,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => readModule1_call_reqs,
      call_acks => readModule1_call_acks,
      return_reqs => readModule1_return_reqs,
      return_acks => readModule1_return_acks,
      call_data  => readModule1_call_data,
      call_tag  => readModule1_call_tag,
      return_tag  => readModule1_return_tag,
      call_mtag => readModule1_tag_in,
      return_mtag => readModule1_tag_out,
      return_data =>readModule1_return_data,
      call_mreq => readModule1_start_req,
      call_mack => readModule1_start_ack,
      return_mreq => readModule1_fin_req,
      return_mack => readModule1_fin_ack,
      call_mdata => readModule1_in_args,
      return_mdata => readModule1_out_args,
      clk => clk, 
      reset => reset --
    ); --
  readModule1_instance:readModule1-- 
    generic map(tag_length => 2)
    port map(-- 
      address => readModule1_address,
      data => readModule1_data,
      start_req => readModule1_start_req,
      start_ack => readModule1_start_ack,
      fin_req => readModule1_fin_req,
      fin_ack => readModule1_fin_ack,
      clk => clk,
      reset => reset,
      memoryModule_call_reqs => memoryModule_call_reqs(0 downto 0),
      memoryModule_call_acks => memoryModule_call_acks(0 downto 0),
      memoryModule_call_data => memoryModule_call_data(96 downto 0),
      memoryModule_call_tag => memoryModule_call_tag(0 downto 0),
      memoryModule_return_reqs => memoryModule_return_reqs(0 downto 0),
      memoryModule_return_acks => memoryModule_return_acks(0 downto 0),
      memoryModule_return_data => memoryModule_return_data(63 downto 0),
      memoryModule_return_tag => memoryModule_return_tag(0 downto 0),
      tag_in => readModule1_tag_in,
      tag_out => readModule1_tag_out-- 
    ); -- 
  -- module readModule_maxPool
  readModule_maxPool_index <= readModule_maxPool_in_args(39 downto 32);
  readModule_maxPool_address <= readModule_maxPool_in_args(31 downto 0);
  readModule_maxPool_out_args <= readModule_maxPool_data ;
  -- call arbiter for module readModule_maxPool
  readModule_maxPool_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 40,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 3--
    )
    port map(-- 
      call_reqs => readModule_maxPool_call_reqs,
      call_acks => readModule_maxPool_call_acks,
      return_reqs => readModule_maxPool_return_reqs,
      return_acks => readModule_maxPool_return_acks,
      call_data  => readModule_maxPool_call_data,
      call_tag  => readModule_maxPool_call_tag,
      return_tag  => readModule_maxPool_return_tag,
      call_mtag => readModule_maxPool_tag_in,
      return_mtag => readModule_maxPool_tag_out,
      return_data =>readModule_maxPool_return_data,
      call_mreq => readModule_maxPool_start_req,
      call_mack => readModule_maxPool_start_ack,
      return_mreq => readModule_maxPool_fin_req,
      return_mack => readModule_maxPool_fin_ack,
      call_mdata => readModule_maxPool_in_args,
      return_mdata => readModule_maxPool_out_args,
      clk => clk, 
      reset => reset --
    ); --
  readModule_maxPool_instance:readModule_maxPool-- 
    generic map(tag_length => 4)
    port map(-- 
      index => readModule_maxPool_index,
      address => readModule_maxPool_address,
      data => readModule_maxPool_data,
      start_req => readModule_maxPool_start_req,
      start_ack => readModule_maxPool_start_ack,
      fin_req => readModule_maxPool_fin_req,
      fin_ack => readModule_maxPool_fin_ack,
      clk => clk,
      reset => reset,
      memoryModule_call_reqs => memoryModule_call_reqs(2 downto 2),
      memoryModule_call_acks => memoryModule_call_acks(2 downto 2),
      memoryModule_call_data => memoryModule_call_data(290 downto 194),
      memoryModule_call_tag => memoryModule_call_tag(2 downto 2),
      memoryModule_return_reqs => memoryModule_return_reqs(2 downto 2),
      memoryModule_return_acks => memoryModule_return_acks(2 downto 2),
      memoryModule_return_data => memoryModule_return_data(191 downto 128),
      memoryModule_return_tag => memoryModule_return_tag(2 downto 2),
      tag_in => readModule_maxPool_tag_in,
      tag_out => readModule_maxPool_tag_out-- 
    ); -- 
  -- module sendOutput
  -- call arbiter for module sendOutput
  sendOutput_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendOutput_call_reqs,
      call_acks => sendOutput_call_acks,
      return_reqs => sendOutput_return_reqs,
      return_acks => sendOutput_return_acks,
      call_tag  => sendOutput_call_tag,
      return_tag  => sendOutput_return_tag,
      call_mtag => sendOutput_tag_in,
      return_mtag => sendOutput_tag_out,
      call_mreq => sendOutput_start_req,
      call_mack => sendOutput_start_ack,
      return_mreq => sendOutput_fin_req,
      return_mack => sendOutput_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  sendOutput_instance:sendOutput-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendOutput_start_req,
      start_ack => sendOutput_start_ack,
      fin_req => sendOutput_fin_req,
      fin_ack => sendOutput_fin_ack,
      clk => clk,
      reset => reset,
      system_output_pipe_pipe_write_req => system_output_pipe_pipe_write_req(1 downto 1),
      system_output_pipe_pipe_write_ack => system_output_pipe_pipe_write_ack(1 downto 1),
      system_output_pipe_pipe_write_data => system_output_pipe_pipe_write_data(15 downto 8),
      readModule1_call_reqs => readModule1_call_reqs(0 downto 0),
      readModule1_call_acks => readModule1_call_acks(0 downto 0),
      readModule1_call_data => readModule1_call_data(31 downto 0),
      readModule1_call_tag => readModule1_call_tag(0 downto 0),
      readModule1_return_reqs => readModule1_return_reqs(0 downto 0),
      readModule1_return_acks => readModule1_return_acks(0 downto 0),
      readModule1_return_data => readModule1_return_data(63 downto 0),
      readModule1_return_tag => readModule1_return_tag(0 downto 0),
      tag_in => sendOutput_tag_in,
      tag_out => sendOutput_tag_out-- 
    ); -- 
  -- module systemTOP
  systemTOP_instance:systemTOP-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => systemTOP_start_req,
      start_ack => systemTOP_start_ack,
      fin_req => systemTOP_fin_req,
      fin_ack => systemTOP_fin_ack,
      clk => clk,
      reset => reset,
      system_output_pipe_pipe_write_req => system_output_pipe_pipe_write_req(0 downto 0),
      system_output_pipe_pipe_write_ack => system_output_pipe_pipe_write_ack(0 downto 0),
      system_output_pipe_pipe_write_data => system_output_pipe_pipe_write_data(7 downto 0),
      fill_input_call_reqs => fill_input_call_reqs(0 downto 0),
      fill_input_call_acks => fill_input_call_acks(0 downto 0),
      fill_input_call_tag => fill_input_call_tag(0 downto 0),
      fill_input_return_reqs => fill_input_return_reqs(0 downto 0),
      fill_input_return_acks => fill_input_return_acks(0 downto 0),
      fill_input_return_tag => fill_input_return_tag(0 downto 0),
      maxPool4_call_reqs => maxPool4_call_reqs(0 downto 0),
      maxPool4_call_acks => maxPool4_call_acks(0 downto 0),
      maxPool4_call_data => maxPool4_call_data(175 downto 0),
      maxPool4_call_tag => maxPool4_call_tag(0 downto 0),
      maxPool4_return_reqs => maxPool4_return_reqs(0 downto 0),
      maxPool4_return_acks => maxPool4_return_acks(0 downto 0),
      maxPool4_return_data => maxPool4_return_data(7 downto 0),
      maxPool4_return_tag => maxPool4_return_tag(0 downto 0),
      sendOutput_call_reqs => sendOutput_call_reqs(0 downto 0),
      sendOutput_call_acks => sendOutput_call_acks(0 downto 0),
      sendOutput_call_tag => sendOutput_call_tag(0 downto 0),
      sendOutput_return_reqs => sendOutput_return_reqs(0 downto 0),
      sendOutput_return_acks => sendOutput_return_acks(0 downto 0),
      sendOutput_return_tag => sendOutput_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => systemTOP_tag_in,
      tag_out => systemTOP_tag_out-- 
    ); -- 
  -- module will be run forever 
  systemTOP_tag_in <= (others => '0');
  systemTOP_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => systemTOP_start_req, start_ack => systemTOP_start_ack,  fin_req => systemTOP_fin_req,  fin_ack => systemTOP_fin_ack);
  -- module timer
  timer_out_args <= timer_T ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      T => timer_T,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      timer_resp_pipe_read_req => timer_resp_pipe_read_req(0 downto 0),
      timer_resp_pipe_read_ack => timer_resp_pipe_read_ack(0 downto 0),
      timer_resp_pipe_read_data => timer_resp_pipe_read_data(63 downto 0),
      timer_req_pipe_write_req => timer_req_pipe_write_req(0 downto 0),
      timer_req_pipe_write_ack => timer_req_pipe_write_ack(0 downto 0),
      timer_req_pipe_write_data => timer_req_pipe_write_data(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      timer_req_pipe_read_req => timer_req_pipe_read_req(0 downto 0),
      timer_req_pipe_read_ack => timer_req_pipe_read_ack(0 downto 0),
      timer_req_pipe_read_data => timer_req_pipe_read_data(0 downto 0),
      timer_resp_pipe_write_req => timer_resp_pipe_write_req(0 downto 0),
      timer_resp_pipe_write_ack => timer_resp_pipe_write_ack(0 downto 0),
      timer_resp_pipe_write_data => timer_resp_pipe_write_data(63 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  -- module writeModule1
  writeModule1_address <= writeModule1_in_args(95 downto 64);
  writeModule1_data <= writeModule1_in_args(63 downto 0);
  -- call arbiter for module writeModule1
  writeModule1_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 96,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writeModule1_call_reqs,
      call_acks => writeModule1_call_acks,
      return_reqs => writeModule1_return_reqs,
      return_acks => writeModule1_return_acks,
      call_data  => writeModule1_call_data,
      call_tag  => writeModule1_call_tag,
      return_tag  => writeModule1_return_tag,
      call_mtag => writeModule1_tag_in,
      return_mtag => writeModule1_tag_out,
      call_mreq => writeModule1_start_req,
      call_mack => writeModule1_start_ack,
      return_mreq => writeModule1_fin_req,
      return_mack => writeModule1_fin_ack,
      call_mdata => writeModule1_in_args,
      clk => clk, 
      reset => reset --
    ); --
  writeModule1_instance:writeModule1-- 
    generic map(tag_length => 2)
    port map(-- 
      address => writeModule1_address,
      data => writeModule1_data,
      start_req => writeModule1_start_req,
      start_ack => writeModule1_start_ack,
      fin_req => writeModule1_fin_req,
      fin_ack => writeModule1_fin_ack,
      clk => clk,
      reset => reset,
      memoryModule_call_reqs => memoryModule_call_reqs(3 downto 3),
      memoryModule_call_acks => memoryModule_call_acks(3 downto 3),
      memoryModule_call_data => memoryModule_call_data(387 downto 291),
      memoryModule_call_tag => memoryModule_call_tag(3 downto 3),
      memoryModule_return_reqs => memoryModule_return_reqs(3 downto 3),
      memoryModule_return_acks => memoryModule_return_acks(3 downto 3),
      memoryModule_return_data => memoryModule_return_data(255 downto 192),
      memoryModule_return_tag => memoryModule_return_tag(3 downto 3),
      tag_in => writeModule1_tag_in,
      tag_out => writeModule1_tag_out-- 
    ); -- 
  -- module writeModule_maxPool
  writeModule_maxPool_index <= writeModule_maxPool_in_args(103 downto 96);
  writeModule_maxPool_address <= writeModule_maxPool_in_args(95 downto 64);
  writeModule_maxPool_data <= writeModule_maxPool_in_args(63 downto 0);
  writeModule_maxPool_out_args <= writeModule_maxPool_done ;
  -- call arbiter for module writeModule_maxPool
  writeModule_maxPool_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 104,
      return_data_width => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writeModule_maxPool_call_reqs,
      call_acks => writeModule_maxPool_call_acks,
      return_reqs => writeModule_maxPool_return_reqs,
      return_acks => writeModule_maxPool_return_acks,
      call_data  => writeModule_maxPool_call_data,
      call_tag  => writeModule_maxPool_call_tag,
      return_tag  => writeModule_maxPool_return_tag,
      call_mtag => writeModule_maxPool_tag_in,
      return_mtag => writeModule_maxPool_tag_out,
      return_data =>writeModule_maxPool_return_data,
      call_mreq => writeModule_maxPool_start_req,
      call_mack => writeModule_maxPool_start_ack,
      return_mreq => writeModule_maxPool_fin_req,
      return_mack => writeModule_maxPool_fin_ack,
      call_mdata => writeModule_maxPool_in_args,
      return_mdata => writeModule_maxPool_out_args,
      clk => clk, 
      reset => reset --
    ); --
  writeModule_maxPool_instance:writeModule_maxPool-- 
    generic map(tag_length => 2)
    port map(-- 
      index => writeModule_maxPool_index,
      address => writeModule_maxPool_address,
      data => writeModule_maxPool_data,
      done => writeModule_maxPool_done,
      start_req => writeModule_maxPool_start_req,
      start_ack => writeModule_maxPool_start_ack,
      fin_req => writeModule_maxPool_fin_req,
      fin_ack => writeModule_maxPool_fin_ack,
      clk => clk,
      reset => reset,
      memoryModule_call_reqs => memoryModule_call_reqs(1 downto 1),
      memoryModule_call_acks => memoryModule_call_acks(1 downto 1),
      memoryModule_call_data => memoryModule_call_data(193 downto 97),
      memoryModule_call_tag => memoryModule_call_tag(1 downto 1),
      memoryModule_return_reqs => memoryModule_return_reqs(1 downto 1),
      memoryModule_return_acks => memoryModule_return_acks(1 downto 1),
      memoryModule_return_data => memoryModule_return_data(127 downto 64),
      memoryModule_return_tag => memoryModule_return_tag(1 downto 1),
      tag_in => writeModule_maxPool_tag_in,
      tag_out => writeModule_maxPool_tag_out-- 
    ); -- 
  MAIN_MEM_REQUEST_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe MAIN_MEM_REQUEST",
      num_reads => 1,
      num_writes => 1,
      data_width => 110,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 16 --
    )
    port map( -- 
      read_req => MAIN_MEM_REQUEST_pipe_read_req,
      read_ack => MAIN_MEM_REQUEST_pipe_read_ack,
      read_data => MAIN_MEM_REQUEST_pipe_read_data,
      write_req => MAIN_MEM_REQUEST_pipe_write_req,
      write_ack => MAIN_MEM_REQUEST_pipe_write_ack,
      write_data => MAIN_MEM_REQUEST_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MAIN_MEM_RESPONSE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe MAIN_MEM_RESPONSE",
      num_reads => 1,
      num_writes => 1,
      data_width => 65,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 16 --
    )
    port map( -- 
      read_req => MAIN_MEM_RESPONSE_pipe_read_req,
      read_ack => MAIN_MEM_RESPONSE_pipe_read_ack,
      read_data => MAIN_MEM_RESPONSE_pipe_read_data,
      write_req => MAIN_MEM_RESPONSE_pipe_write_req,
      write_ack => MAIN_MEM_RESPONSE_pipe_write_ack,
      write_data => MAIN_MEM_RESPONSE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  system_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe system_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => system_input_pipe_pipe_read_req,
      read_ack => system_input_pipe_pipe_read_ack,
      read_data => system_input_pipe_pipe_read_data,
      write_req => system_input_pipe_pipe_write_req,
      write_ack => system_input_pipe_pipe_write_ack,
      write_data => system_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  system_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe system_output_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => system_output_pipe_pipe_read_req,
      read_ack => system_output_pipe_pipe_read_ack,
      read_data => system_output_pipe_pipe_read_data,
      write_req => system_output_pipe_pipe_write_req,
      write_ack => system_output_pipe_pipe_write_ack,
      write_data => system_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  timer_req_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_req",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_req_pipe_read_req,
      read_ack => timer_req_pipe_read_ack,
      read_data => timer_req_pipe_read_data,
      write_req => timer_req_pipe_write_req,
      write_ack => timer_req_pipe_write_ack,
      write_data => timer_req_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  timer_resp_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_resp",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_resp_pipe_read_req,
      read_ack => timer_resp_pipe_read_ack,
      read_data => timer_resp_pipe_read_data,
      write_req => timer_resp_pipe_write_req,
      write_ack => timer_resp_pipe_write_ack,
      write_data => timer_resp_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  -- 
end ahir_system_arch;
