-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_39_start: Boolean;
  signal convTranspose_CP_39_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal addr_of_538_final_reg_ack_0 : boolean;
  signal addr_of_538_final_reg_req_0 : boolean;
  signal type_cast_548_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_872_inst_req_0 : boolean;
  signal type_cast_374_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_543_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_543_inst_ack_1 : boolean;
  signal type_cast_390_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_872_inst_ack_1 : boolean;
  signal addr_of_538_final_reg_ack_1 : boolean;
  signal type_cast_837_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_895_inst_req_0 : boolean;
  signal type_cast_390_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_354_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_895_inst_ack_0 : boolean;
  signal array_obj_ref_1302_index_offset_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_352_inst_req_0 : boolean;
  signal type_cast_374_inst_req_1 : boolean;
  signal type_cast_1007_inst_req_1 : boolean;
  signal type_cast_452_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_851_inst_req_0 : boolean;
  signal type_cast_1235_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_543_inst_ack_0 : boolean;
  signal type_cast_548_inst_ack_0 : boolean;
  signal type_cast_548_inst_req_1 : boolean;
  signal type_cast_548_inst_ack_1 : boolean;
  signal type_cast_900_inst_req_0 : boolean;
  signal type_cast_958_inst_ack_0 : boolean;
  signal type_cast_816_inst_req_0 : boolean;
  signal type_cast_42_inst_req_0 : boolean;
  signal type_cast_921_inst_req_1 : boolean;
  signal type_cast_452_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_914_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_383_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_383_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_383_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_383_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_352_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_352_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_352_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_req_0 : boolean;
  signal type_cast_405_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_ack_1 : boolean;
  signal addr_of_538_final_reg_req_1 : boolean;
  signal array_obj_ref_1036_index_offset_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_37_inst_req_0 : boolean;
  signal type_cast_405_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_37_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_37_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_37_inst_ack_1 : boolean;
  signal type_cast_954_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_115_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_115_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_369_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_115_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_115_inst_ack_1 : boolean;
  signal if_stmt_481_branch_ack_1 : boolean;
  signal type_cast_42_inst_ack_0 : boolean;
  signal type_cast_42_inst_req_1 : boolean;
  signal type_cast_42_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_851_inst_req_1 : boolean;
  signal type_cast_374_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_51_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_51_inst_ack_0 : boolean;
  signal type_cast_374_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_51_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_51_inst_ack_1 : boolean;
  signal type_cast_508_inst_ack_1 : boolean;
  signal type_cast_508_inst_req_1 : boolean;
  signal type_cast_452_inst_ack_0 : boolean;
  signal type_cast_958_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_53_inst_req_0 : boolean;
  signal type_cast_405_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_53_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_53_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_53_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_369_inst_ack_1 : boolean;
  signal type_cast_958_inst_req_1 : boolean;
  signal type_cast_58_inst_req_0 : boolean;
  signal type_cast_405_inst_req_0 : boolean;
  signal type_cast_58_inst_ack_0 : boolean;
  signal type_cast_58_inst_req_1 : boolean;
  signal type_cast_58_inst_ack_1 : boolean;
  signal type_cast_816_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_66_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_66_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_66_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_66_inst_ack_1 : boolean;
  signal type_cast_508_inst_ack_0 : boolean;
  signal type_cast_508_inst_req_0 : boolean;
  signal type_cast_452_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_431_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_68_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_68_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_68_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_68_inst_ack_1 : boolean;
  signal type_cast_900_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1196_inst_req_1 : boolean;
  signal type_cast_73_inst_req_0 : boolean;
  signal type_cast_73_inst_ack_0 : boolean;
  signal type_cast_73_inst_req_1 : boolean;
  signal type_cast_73_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1227_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_431_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_82_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_82_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_82_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_82_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_84_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_84_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_84_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_84_inst_ack_1 : boolean;
  signal addr_of_1303_final_reg_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_445_inst_ack_1 : boolean;
  signal type_cast_89_inst_req_0 : boolean;
  signal type_cast_89_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_445_inst_req_1 : boolean;
  signal type_cast_89_inst_req_1 : boolean;
  signal type_cast_89_inst_ack_1 : boolean;
  signal ptr_deref_929_store_0_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_369_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_431_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_431_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_ack_1 : boolean;
  signal addr_of_1037_final_reg_req_0 : boolean;
  signal addr_of_1303_final_reg_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_99_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_99_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_99_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_99_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_853_inst_req_1 : boolean;
  signal type_cast_104_inst_req_0 : boolean;
  signal type_cast_104_inst_ack_0 : boolean;
  signal type_cast_104_inst_req_1 : boolean;
  signal type_cast_104_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_416_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_113_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_113_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_369_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_113_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_113_inst_ack_1 : boolean;
  signal if_stmt_481_branch_ack_0 : boolean;
  signal type_cast_436_inst_ack_1 : boolean;
  signal type_cast_261_inst_req_0 : boolean;
  signal type_cast_261_inst_ack_0 : boolean;
  signal type_cast_261_inst_req_1 : boolean;
  signal type_cast_261_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_872_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_830_inst_ack_0 : boolean;
  signal type_cast_436_inst_req_1 : boolean;
  signal type_cast_275_inst_req_0 : boolean;
  signal type_cast_275_inst_ack_0 : boolean;
  signal type_cast_275_inst_req_1 : boolean;
  signal type_cast_275_inst_ack_1 : boolean;
  signal type_cast_954_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_914_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_416_inst_req_1 : boolean;
  signal type_cast_120_inst_req_0 : boolean;
  signal type_cast_120_inst_ack_0 : boolean;
  signal type_cast_120_inst_req_1 : boolean;
  signal type_cast_120_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1208_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_130_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_130_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_130_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_400_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_130_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_830_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_874_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_445_inst_ack_0 : boolean;
  signal type_cast_135_inst_req_0 : boolean;
  signal type_cast_135_inst_ack_0 : boolean;
  signal type_cast_135_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_400_inst_req_1 : boolean;
  signal type_cast_135_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_416_inst_ack_0 : boolean;
  signal type_cast_921_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_144_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_144_inst_ack_0 : boolean;
  signal type_cast_962_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_144_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_144_inst_ack_1 : boolean;
  signal if_stmt_481_branch_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_146_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_146_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_146_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_146_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_811_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_914_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_416_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_445_inst_req_0 : boolean;
  signal type_cast_151_inst_req_0 : boolean;
  signal type_cast_151_inst_ack_0 : boolean;
  signal type_cast_151_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_400_inst_ack_0 : boolean;
  signal type_cast_151_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_541_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_429_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_367_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_400_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_429_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_161_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_161_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_367_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_161_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_161_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_895_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_385_inst_ack_1 : boolean;
  signal type_cast_166_inst_req_0 : boolean;
  signal type_cast_166_inst_ack_0 : boolean;
  signal type_cast_166_inst_req_1 : boolean;
  signal type_cast_166_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_541_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_175_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_175_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_175_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_175_inst_ack_1 : boolean;
  signal type_cast_1007_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_429_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_429_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_177_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_177_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_367_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_177_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_177_inst_ack_1 : boolean;
  signal array_obj_ref_537_index_offset_ack_1 : boolean;
  signal type_cast_182_inst_req_0 : boolean;
  signal type_cast_182_inst_ack_0 : boolean;
  signal type_cast_182_inst_req_1 : boolean;
  signal type_cast_182_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_367_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_190_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_190_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_190_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_190_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_916_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1227_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_447_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_874_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_192_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_192_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_192_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_192_inst_ack_1 : boolean;
  signal array_obj_ref_537_index_offset_req_1 : boolean;
  signal if_stmt_466_branch_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_853_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_385_inst_req_1 : boolean;
  signal type_cast_958_inst_ack_1 : boolean;
  signal type_cast_197_inst_req_0 : boolean;
  signal type_cast_197_inst_ack_0 : boolean;
  signal type_cast_197_inst_req_1 : boolean;
  signal type_cast_197_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_206_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_206_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_206_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_206_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_916_inst_ack_1 : boolean;
  signal if_stmt_466_branch_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_447_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_830_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_208_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_208_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_208_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_208_inst_ack_1 : boolean;
  signal type_cast_900_inst_req_1 : boolean;
  signal type_cast_213_inst_req_0 : boolean;
  signal type_cast_213_inst_ack_0 : boolean;
  signal type_cast_213_inst_req_1 : boolean;
  signal type_cast_858_inst_req_0 : boolean;
  signal type_cast_213_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_541_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_853_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_221_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_221_inst_ack_0 : boolean;
  signal type_cast_359_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_221_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_221_inst_ack_1 : boolean;
  signal array_obj_ref_1036_index_offset_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_447_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_223_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_398_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_223_inst_ack_0 : boolean;
  signal type_cast_359_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_223_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_223_inst_ack_1 : boolean;
  signal array_obj_ref_537_index_offset_ack_0 : boolean;
  signal if_stmt_466_branch_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_872_inst_ack_0 : boolean;
  signal type_cast_900_inst_ack_1 : boolean;
  signal type_cast_228_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_398_inst_req_1 : boolean;
  signal type_cast_228_inst_ack_0 : boolean;
  signal type_cast_228_inst_req_1 : boolean;
  signal type_cast_858_inst_ack_0 : boolean;
  signal type_cast_228_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_541_inst_req_0 : boolean;
  signal type_cast_421_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_237_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_237_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_237_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_237_inst_ack_1 : boolean;
  signal array_obj_ref_537_index_offset_req_0 : boolean;
  signal type_cast_954_inst_req_1 : boolean;
  signal type_cast_816_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_447_inst_req_0 : boolean;
  signal type_cast_421_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_239_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_239_inst_ack_0 : boolean;
  signal type_cast_359_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_239_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_398_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_239_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_414_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_385_inst_ack_0 : boolean;
  signal type_cast_244_inst_req_0 : boolean;
  signal type_cast_244_inst_ack_0 : boolean;
  signal type_cast_244_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_398_inst_req_0 : boolean;
  signal type_cast_244_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_851_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_414_inst_req_1 : boolean;
  signal type_cast_253_inst_req_0 : boolean;
  signal type_cast_253_inst_ack_0 : boolean;
  signal type_cast_253_inst_req_1 : boolean;
  signal type_cast_359_inst_req_0 : boolean;
  signal type_cast_253_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_414_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_414_inst_req_0 : boolean;
  signal type_cast_257_inst_req_0 : boolean;
  signal type_cast_257_inst_ack_0 : boolean;
  signal type_cast_257_inst_req_1 : boolean;
  signal type_cast_257_inst_ack_1 : boolean;
  signal type_cast_436_inst_ack_0 : boolean;
  signal type_cast_279_inst_req_0 : boolean;
  signal type_cast_279_inst_ack_0 : boolean;
  signal type_cast_279_inst_req_1 : boolean;
  signal type_cast_279_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_543_inst_req_0 : boolean;
  signal ptr_deref_929_store_0_req_1 : boolean;
  signal type_cast_436_inst_req_0 : boolean;
  signal type_cast_283_inst_req_0 : boolean;
  signal type_cast_283_inst_ack_0 : boolean;
  signal type_cast_283_inst_req_1 : boolean;
  signal type_cast_283_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_385_inst_req_0 : boolean;
  signal if_stmt_943_branch_req_0 : boolean;
  signal type_cast_1273_inst_ack_1 : boolean;
  signal type_cast_287_inst_req_0 : boolean;
  signal type_cast_287_inst_ack_0 : boolean;
  signal type_cast_858_inst_req_1 : boolean;
  signal type_cast_287_inst_req_1 : boolean;
  signal type_cast_287_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_305_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_305_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_305_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_305_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_895_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_851_inst_ack_1 : boolean;
  signal type_cast_421_inst_ack_0 : boolean;
  signal type_cast_421_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_307_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_307_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_307_inst_req_1 : boolean;
  signal type_cast_390_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_307_inst_ack_1 : boolean;
  signal type_cast_962_inst_req_1 : boolean;
  signal type_cast_921_inst_req_0 : boolean;
  signal type_cast_312_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_914_inst_req_0 : boolean;
  signal type_cast_312_inst_ack_0 : boolean;
  signal type_cast_312_inst_req_1 : boolean;
  signal type_cast_390_inst_req_1 : boolean;
  signal type_cast_312_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_354_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_354_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_321_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_321_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_321_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_321_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_323_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_323_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_323_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_323_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_354_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_853_inst_req_0 : boolean;
  signal type_cast_328_inst_req_0 : boolean;
  signal type_cast_328_inst_ack_0 : boolean;
  signal type_cast_328_inst_req_1 : boolean;
  signal type_cast_328_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_830_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_336_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_336_inst_ack_0 : boolean;
  signal type_cast_858_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_336_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_336_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1196_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_338_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_338_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_338_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_338_inst_ack_1 : boolean;
  signal type_cast_343_inst_req_0 : boolean;
  signal type_cast_343_inst_ack_0 : boolean;
  signal type_cast_343_inst_req_1 : boolean;
  signal type_cast_343_inst_ack_1 : boolean;
  signal type_cast_954_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_557_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_557_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_557_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_557_inst_ack_1 : boolean;
  signal array_obj_ref_1036_index_offset_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_559_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_559_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_559_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_559_inst_ack_1 : boolean;
  signal array_obj_ref_1036_index_offset_req_0 : boolean;
  signal type_cast_962_inst_ack_0 : boolean;
  signal type_cast_564_inst_req_0 : boolean;
  signal type_cast_564_inst_ack_0 : boolean;
  signal type_cast_564_inst_req_1 : boolean;
  signal type_cast_564_inst_ack_1 : boolean;
  signal array_obj_ref_1302_index_offset_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_578_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_578_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_578_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_578_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1211_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_580_inst_req_0 : boolean;
  signal ptr_deref_929_store_0_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_580_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_580_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_580_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1196_inst_req_0 : boolean;
  signal type_cast_962_inst_req_0 : boolean;
  signal type_cast_585_inst_req_0 : boolean;
  signal ptr_deref_929_store_0_req_0 : boolean;
  signal type_cast_585_inst_ack_0 : boolean;
  signal type_cast_585_inst_req_1 : boolean;
  signal type_cast_585_inst_ack_1 : boolean;
  signal array_obj_ref_1302_index_offset_ack_0 : boolean;
  signal type_cast_837_inst_req_1 : boolean;
  signal addr_of_1303_final_reg_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_599_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_599_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_599_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_599_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1211_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_601_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_601_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_601_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_601_inst_ack_1 : boolean;
  signal if_stmt_980_branch_ack_0 : boolean;
  signal type_cast_606_inst_req_0 : boolean;
  signal type_cast_606_inst_ack_0 : boolean;
  signal type_cast_606_inst_req_1 : boolean;
  signal type_cast_606_inst_ack_1 : boolean;
  signal type_cast_1007_inst_ack_0 : boolean;
  signal type_cast_837_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_620_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_620_inst_ack_0 : boolean;
  signal type_cast_837_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_620_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_620_inst_ack_1 : boolean;
  signal addr_of_1037_final_reg_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_622_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_622_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_622_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_622_inst_ack_1 : boolean;
  signal addr_of_1037_final_reg_req_1 : boolean;
  signal addr_of_1303_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_893_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_893_inst_req_1 : boolean;
  signal type_cast_627_inst_req_0 : boolean;
  signal type_cast_627_inst_ack_0 : boolean;
  signal type_cast_627_inst_req_1 : boolean;
  signal type_cast_627_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1227_inst_req_1 : boolean;
  signal if_stmt_943_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_641_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_641_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_641_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_641_inst_ack_1 : boolean;
  signal if_stmt_980_branch_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_643_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_643_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_643_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_643_inst_ack_1 : boolean;
  signal type_cast_1235_inst_req_0 : boolean;
  signal RPIPE_Block3_done_1227_inst_ack_1 : boolean;
  signal type_cast_648_inst_req_0 : boolean;
  signal type_cast_648_inst_ack_0 : boolean;
  signal type_cast_648_inst_req_1 : boolean;
  signal type_cast_648_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_893_inst_ack_0 : boolean;
  signal type_cast_1007_inst_req_0 : boolean;
  signal array_obj_ref_1302_index_offset_req_1 : boolean;
  signal addr_of_1037_final_reg_ack_0 : boolean;
  signal if_stmt_943_branch_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_662_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_662_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_662_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_662_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_664_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_664_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_664_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_664_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_893_inst_req_0 : boolean;
  signal type_cast_669_inst_req_0 : boolean;
  signal type_cast_669_inst_ack_0 : boolean;
  signal type_cast_669_inst_req_1 : boolean;
  signal type_cast_669_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_832_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1208_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_683_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_683_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_832_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_683_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_683_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_685_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_685_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_685_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_685_inst_ack_1 : boolean;
  signal if_stmt_980_branch_req_0 : boolean;
  signal type_cast_690_inst_req_0 : boolean;
  signal type_cast_690_inst_ack_0 : boolean;
  signal type_cast_690_inst_req_1 : boolean;
  signal type_cast_690_inst_ack_1 : boolean;
  signal type_cast_879_inst_ack_1 : boolean;
  signal type_cast_879_inst_req_1 : boolean;
  signal type_cast_921_inst_ack_1 : boolean;
  signal ptr_deref_698_store_0_req_0 : boolean;
  signal ptr_deref_698_store_0_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_811_inst_req_1 : boolean;
  signal type_cast_816_inst_ack_0 : boolean;
  signal ptr_deref_698_store_0_req_1 : boolean;
  signal type_cast_879_inst_ack_0 : boolean;
  signal ptr_deref_698_store_0_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_832_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_832_inst_req_0 : boolean;
  signal type_cast_879_inst_req_0 : boolean;
  signal type_cast_1273_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1196_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_874_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_874_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_916_inst_ack_0 : boolean;
  signal if_stmt_712_branch_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_916_inst_req_0 : boolean;
  signal if_stmt_712_branch_ack_1 : boolean;
  signal if_stmt_712_branch_ack_0 : boolean;
  signal type_cast_1235_inst_req_1 : boolean;
  signal type_cast_739_inst_req_0 : boolean;
  signal type_cast_739_inst_ack_0 : boolean;
  signal type_cast_739_inst_req_1 : boolean;
  signal type_cast_739_inst_ack_1 : boolean;
  signal call_stmt_1231_call_req_0 : boolean;
  signal WPIPE_Block3_start_1208_inst_req_1 : boolean;
  signal call_stmt_1231_call_ack_0 : boolean;
  signal type_cast_1235_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1208_inst_ack_1 : boolean;
  signal array_obj_ref_768_index_offset_req_0 : boolean;
  signal array_obj_ref_768_index_offset_ack_0 : boolean;
  signal array_obj_ref_768_index_offset_req_1 : boolean;
  signal array_obj_ref_768_index_offset_ack_1 : boolean;
  signal addr_of_769_final_reg_req_0 : boolean;
  signal addr_of_769_final_reg_ack_0 : boolean;
  signal addr_of_769_final_reg_req_1 : boolean;
  signal addr_of_769_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_772_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_772_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_772_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_772_inst_ack_1 : boolean;
  signal call_stmt_1231_call_req_1 : boolean;
  signal call_stmt_1231_call_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_774_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_774_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1211_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_774_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_774_inst_ack_1 : boolean;
  signal type_cast_779_inst_req_0 : boolean;
  signal type_cast_779_inst_ack_0 : boolean;
  signal type_cast_779_inst_req_1 : boolean;
  signal type_cast_779_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_788_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_788_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_788_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_788_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_790_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_790_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_790_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_790_inst_ack_1 : boolean;
  signal type_cast_795_inst_req_0 : boolean;
  signal type_cast_795_inst_ack_0 : boolean;
  signal type_cast_795_inst_req_1 : boolean;
  signal type_cast_795_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_809_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_809_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_809_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_809_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_811_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_811_inst_ack_0 : boolean;
  signal RPIPE_Block2_done_1224_inst_ack_1 : boolean;
  signal RPIPE_Block2_done_1224_inst_req_1 : boolean;
  signal type_cast_1273_inst_ack_0 : boolean;
  signal type_cast_1273_inst_req_0 : boolean;
  signal ptr_deref_1040_store_0_req_0 : boolean;
  signal RPIPE_Block2_done_1224_inst_ack_0 : boolean;
  signal ptr_deref_1040_store_0_ack_0 : boolean;
  signal WPIPE_Block3_start_1193_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1211_inst_ack_0 : boolean;
  signal ptr_deref_1040_store_0_req_1 : boolean;
  signal RPIPE_Block2_done_1224_inst_req_0 : boolean;
  signal ptr_deref_1040_store_0_ack_1 : boolean;
  signal WPIPE_Block3_start_1205_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1205_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1193_inst_req_1 : boolean;
  signal if_stmt_1055_branch_req_0 : boolean;
  signal if_stmt_1055_branch_ack_1 : boolean;
  signal if_stmt_1055_branch_ack_0 : boolean;
  signal call_stmt_1066_call_req_0 : boolean;
  signal call_stmt_1066_call_ack_0 : boolean;
  signal call_stmt_1066_call_req_1 : boolean;
  signal call_stmt_1066_call_ack_1 : boolean;
  signal WPIPE_Block3_start_1205_inst_ack_0 : boolean;
  signal type_cast_1071_inst_req_0 : boolean;
  signal type_cast_1071_inst_ack_0 : boolean;
  signal type_cast_1071_inst_req_1 : boolean;
  signal type_cast_1071_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1205_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1073_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1073_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1073_inst_req_1 : boolean;
  signal if_stmt_1246_branch_ack_0 : boolean;
  signal WPIPE_Block0_start_1073_inst_ack_1 : boolean;
  signal RPIPE_Block1_done_1221_inst_ack_1 : boolean;
  signal RPIPE_Block1_done_1221_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1076_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1076_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1076_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1076_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1079_inst_req_0 : boolean;
  signal if_stmt_1246_branch_ack_1 : boolean;
  signal WPIPE_Block0_start_1079_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1079_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1079_inst_ack_1 : boolean;
  signal ptr_deref_1307_load_0_ack_1 : boolean;
  signal ptr_deref_1307_load_0_req_1 : boolean;
  signal RPIPE_Block1_done_1221_inst_ack_0 : boolean;
  signal RPIPE_Block1_done_1221_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1082_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1082_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1202_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1082_inst_req_1 : boolean;
  signal if_stmt_1246_branch_req_0 : boolean;
  signal WPIPE_Block0_start_1082_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1202_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1085_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1085_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1085_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1085_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1088_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1088_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1202_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1088_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1088_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1202_inst_req_0 : boolean;
  signal ptr_deref_1307_load_0_ack_0 : boolean;
  signal ptr_deref_1307_load_0_req_0 : boolean;
  signal RPIPE_Block0_done_1218_inst_ack_1 : boolean;
  signal RPIPE_Block0_done_1218_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1091_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1091_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1091_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1242_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1091_inst_ack_1 : boolean;
  signal RPIPE_Block0_done_1218_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1094_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1242_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1094_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1094_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1094_inst_ack_1 : boolean;
  signal RPIPE_Block0_done_1218_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1097_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1097_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1097_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1242_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1097_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1100_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1242_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1100_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1100_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1100_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1199_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1214_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1214_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1103_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1103_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1199_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1103_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1103_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1214_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1106_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1106_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1106_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1106_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1199_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1214_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1109_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1109_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1199_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1109_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1109_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1112_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1112_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1112_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1112_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1115_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1115_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1115_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1115_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1118_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1118_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1118_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1118_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1121_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1121_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1121_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1121_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1124_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1124_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1124_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1124_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1127_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1127_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1127_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1127_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1130_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1130_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1130_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1130_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1133_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1133_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1133_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1133_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1136_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1136_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1136_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1136_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1139_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1139_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1139_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1139_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1142_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1142_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1142_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1142_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1145_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1145_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1145_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1145_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1148_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1148_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1148_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1148_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1151_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1151_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1151_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1151_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1154_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1154_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1154_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1154_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1157_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1157_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1157_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1157_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1160_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1160_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1160_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1160_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1163_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1163_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1163_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1163_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1166_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1166_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1166_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1166_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1169_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1169_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1169_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1169_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1172_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1172_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1172_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1172_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1175_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1175_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1175_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1175_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1178_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1178_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1178_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1178_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1181_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1181_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1181_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1181_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1184_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1184_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1184_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1184_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1187_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1187_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1187_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1187_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1190_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1190_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1190_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1190_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1193_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1193_inst_ack_0 : boolean;
  signal type_cast_1311_inst_req_0 : boolean;
  signal type_cast_1311_inst_ack_0 : boolean;
  signal type_cast_1311_inst_req_1 : boolean;
  signal type_cast_1311_inst_ack_1 : boolean;
  signal type_cast_1321_inst_req_0 : boolean;
  signal type_cast_1321_inst_ack_0 : boolean;
  signal type_cast_1321_inst_req_1 : boolean;
  signal type_cast_1321_inst_ack_1 : boolean;
  signal type_cast_1331_inst_req_0 : boolean;
  signal type_cast_1331_inst_ack_0 : boolean;
  signal type_cast_1331_inst_req_1 : boolean;
  signal type_cast_1331_inst_ack_1 : boolean;
  signal type_cast_1341_inst_req_0 : boolean;
  signal type_cast_1341_inst_ack_0 : boolean;
  signal type_cast_1341_inst_req_1 : boolean;
  signal type_cast_1341_inst_ack_1 : boolean;
  signal type_cast_1351_inst_req_0 : boolean;
  signal type_cast_1351_inst_ack_0 : boolean;
  signal type_cast_1351_inst_req_1 : boolean;
  signal type_cast_1351_inst_ack_1 : boolean;
  signal type_cast_1361_inst_req_0 : boolean;
  signal type_cast_1361_inst_ack_0 : boolean;
  signal type_cast_1361_inst_req_1 : boolean;
  signal type_cast_1361_inst_ack_1 : boolean;
  signal type_cast_1371_inst_req_0 : boolean;
  signal type_cast_1371_inst_ack_0 : boolean;
  signal type_cast_1371_inst_req_1 : boolean;
  signal type_cast_1371_inst_ack_1 : boolean;
  signal type_cast_1381_inst_req_0 : boolean;
  signal type_cast_1381_inst_ack_0 : boolean;
  signal type_cast_1381_inst_req_1 : boolean;
  signal type_cast_1381_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1383_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1383_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1383_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1383_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1386_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1386_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1386_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1386_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1389_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1389_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1389_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1389_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1392_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1392_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1392_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1392_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1395_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1395_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1395_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1395_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1398_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1398_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1398_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1398_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1401_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1401_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1401_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1401_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1404_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1404_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1404_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1404_inst_ack_1 : boolean;
  signal if_stmt_1418_branch_req_0 : boolean;
  signal if_stmt_1418_branch_ack_1 : boolean;
  signal if_stmt_1418_branch_ack_0 : boolean;
  signal phi_stmt_525_req_0 : boolean;
  signal type_cast_531_inst_req_0 : boolean;
  signal type_cast_531_inst_ack_0 : boolean;
  signal type_cast_531_inst_req_1 : boolean;
  signal type_cast_531_inst_ack_1 : boolean;
  signal phi_stmt_525_req_1 : boolean;
  signal phi_stmt_525_ack_0 : boolean;
  signal phi_stmt_756_req_0 : boolean;
  signal type_cast_762_inst_req_0 : boolean;
  signal type_cast_762_inst_ack_0 : boolean;
  signal type_cast_762_inst_req_1 : boolean;
  signal type_cast_762_inst_ack_1 : boolean;
  signal phi_stmt_756_req_1 : boolean;
  signal phi_stmt_756_ack_0 : boolean;
  signal phi_stmt_1024_req_0 : boolean;
  signal type_cast_1030_inst_req_0 : boolean;
  signal type_cast_1030_inst_ack_0 : boolean;
  signal type_cast_1030_inst_req_1 : boolean;
  signal type_cast_1030_inst_ack_1 : boolean;
  signal phi_stmt_1024_req_1 : boolean;
  signal phi_stmt_1024_ack_0 : boolean;
  signal phi_stmt_1290_req_1 : boolean;
  signal type_cast_1293_inst_req_0 : boolean;
  signal type_cast_1293_inst_ack_0 : boolean;
  signal type_cast_1293_inst_req_1 : boolean;
  signal type_cast_1293_inst_ack_1 : boolean;
  signal phi_stmt_1290_req_0 : boolean;
  signal phi_stmt_1290_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_39_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_39: Block -- control-path 
    signal convTranspose_CP_39_elements: BooleanArray(542 downto 0);
    -- 
  begin -- 
    convTranspose_CP_39_elements(0) <= convTranspose_CP_39_start;
    convTranspose_CP_39_symbol <= convTranspose_CP_39_elements(542);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	27 
    -- CP-element group 0: 	34 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	41 
    -- CP-element group 0: 	55 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	153 
    -- CP-element group 0: 	160 
    -- CP-element group 0: 	167 
    -- CP-element group 0: 	174 
    -- CP-element group 0: 	181 
    -- CP-element group 0: 	188 
    -- CP-element group 0: 	90 
    -- CP-element group 0: 	69 
    -- CP-element group 0: 	76 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	100 
    -- CP-element group 0: 	62 
    -- CP-element group 0: 	146 
    -- CP-element group 0: 	139 
    -- CP-element group 0: 	83 
    -- CP-element group 0: 	112 
    -- CP-element group 0: 	115 
    -- CP-element group 0: 	118 
    -- CP-element group 0: 	103 
    -- CP-element group 0: 	106 
    -- CP-element group 0: 	109 
    -- CP-element group 0: 	132 
    -- CP-element group 0: 	125 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	13 
    -- CP-element group 0:  members (101) 
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_390_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_374_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_42_update_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_33/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/branch_block_stmt_33__entry__
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_452_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465__entry__
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_35_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_35_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_35_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_421_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_452_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_405_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_374_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_42_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_42_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_405_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_58_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_58_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_58_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_374_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_73_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_73_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_73_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_405_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_89_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_89_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_89_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_452_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_104_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_104_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_104_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_261_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_261_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_275_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_436_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_275_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_436_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_275_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_120_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_120_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_120_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_135_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_135_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_135_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_253_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_151_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_151_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_151_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_166_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_166_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_166_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_182_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_182_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_182_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_197_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_197_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_197_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_213_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_213_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_213_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_359_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_228_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_228_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_228_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_359_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_421_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_244_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_244_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_244_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_253_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_253_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_257_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_257_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_257_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_261_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_279_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_279_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_279_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_283_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_283_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_283_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_287_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_287_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_287_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_421_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_359_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_312_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_312_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_436_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_312_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_390_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_390_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_328_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_328_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_328_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_343_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_343_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_343_Update/cr
      -- 
    cr_1020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_374_inst_req_1); -- 
    cr_1230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_452_inst_req_1); -- 
    rr_133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => RPIPE_ConvTranspose_input_pipe_35_inst_req_0); -- 
    cr_1104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_405_inst_req_1); -- 
    cr_166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_42_inst_req_1); -- 
    cr_208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_58_inst_req_1); -- 
    cr_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_73_inst_req_1); -- 
    cr_292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_89_inst_req_1); -- 
    cr_334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_104_inst_req_1); -- 
    cr_754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_261_inst_req_1); -- 
    cr_1188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_436_inst_req_1); -- 
    cr_768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_275_inst_req_1); -- 
    cr_376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_120_inst_req_1); -- 
    cr_418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_135_inst_req_1); -- 
    cr_460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_151_inst_req_1); -- 
    cr_502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_166_inst_req_1); -- 
    cr_544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_182_inst_req_1); -- 
    cr_586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_197_inst_req_1); -- 
    cr_628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_213_inst_req_1); -- 
    cr_978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_359_inst_req_1); -- 
    cr_670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_228_inst_req_1); -- 
    cr_1146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_421_inst_req_1); -- 
    cr_712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_244_inst_req_1); -- 
    cr_726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_253_inst_req_1); -- 
    cr_740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_257_inst_req_1); -- 
    cr_782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_279_inst_req_1); -- 
    cr_796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_283_inst_req_1); -- 
    cr_810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_287_inst_req_1); -- 
    cr_852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_312_inst_req_1); -- 
    cr_1062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_390_inst_req_1); -- 
    cr_894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_328_inst_req_1); -- 
    cr_936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_343_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_35_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_35_update_start_
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_35_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_35_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_35_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_35_Update/cr
      -- 
    ra_134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_35_inst_ack_0, ack => convTranspose_CP_39_elements(1)); -- 
    cr_138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(1), ack => RPIPE_ConvTranspose_input_pipe_35_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	7 
    -- CP-element group 2:  members (12) 
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_42_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_42_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_42_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_35_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_35_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_35_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_37_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_37_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_37_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_51_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_51_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_51_Sample/rr
      -- 
    ca_139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_35_inst_ack_1, ack => convTranspose_CP_39_elements(2)); -- 
    req_147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => WPIPE_ConvTranspose_output_pipe_37_inst_req_0); -- 
    rr_161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => type_cast_42_inst_req_0); -- 
    rr_175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => RPIPE_ConvTranspose_input_pipe_51_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_37_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_37_update_start_
      -- CP-element group 3: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_37_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_37_Sample/ack
      -- CP-element group 3: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_37_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_37_Update/req
      -- 
    ack_148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_37_inst_ack_0, ack => convTranspose_CP_39_elements(3)); -- 
    req_152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(3), ack => WPIPE_ConvTranspose_output_pipe_37_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	9 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_37_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_37_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_37_Update/ack
      -- 
    ack_153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_37_inst_ack_1, ack => convTranspose_CP_39_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_42_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_42_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_42_Sample/ra
      -- 
    ra_162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_42_inst_ack_0, ack => convTranspose_CP_39_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	98 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_42_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_42_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_42_Update/ca
      -- 
    ca_167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_42_inst_ack_1, ack => convTranspose_CP_39_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_51_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_51_update_start_
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_51_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_51_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_51_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_51_Update/cr
      -- 
    ra_176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_51_inst_ack_0, ack => convTranspose_CP_39_elements(7)); -- 
    cr_180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(7), ack => RPIPE_ConvTranspose_input_pipe_51_inst_req_1); -- 
    -- CP-element group 8:  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: 	12 
    -- CP-element group 8: 	14 
    -- CP-element group 8:  members (9) 
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_51_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_51_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_51_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_58_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_58_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_58_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_66_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_66_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_66_Sample/rr
      -- 
    ca_181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_51_inst_ack_1, ack => convTranspose_CP_39_elements(8)); -- 
    rr_203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(8), ack => type_cast_58_inst_req_0); -- 
    rr_217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(8), ack => RPIPE_ConvTranspose_input_pipe_66_inst_req_0); -- 
    -- CP-element group 9:  join  transition  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	4 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_53_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_53_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_53_Sample/req
      -- 
    req_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(9), ack => WPIPE_ConvTranspose_output_pipe_53_inst_req_0); -- 
    convTranspose_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "convTranspose_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(4) & convTranspose_CP_39_elements(8);
      gj_convTranspose_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_53_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_53_update_start_
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_53_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_53_Sample/ack
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_53_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_53_Update/req
      -- 
    ack_190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_53_inst_ack_0, ack => convTranspose_CP_39_elements(10)); -- 
    req_194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(10), ack => WPIPE_ConvTranspose_output_pipe_53_inst_req_1); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	16 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_53_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_53_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_53_Update/ack
      -- 
    ack_195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_53_inst_ack_1, ack => convTranspose_CP_39_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	8 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_58_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_58_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_58_Sample/ra
      -- 
    ra_204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_58_inst_ack_0, ack => convTranspose_CP_39_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	98 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_58_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_58_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_58_Update/ca
      -- 
    ca_209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_58_inst_ack_1, ack => convTranspose_CP_39_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	8 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_66_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_66_update_start_
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_66_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_66_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_66_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_66_Update/cr
      -- 
    ra_218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_66_inst_ack_0, ack => convTranspose_CP_39_elements(14)); -- 
    cr_222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(14), ack => RPIPE_ConvTranspose_input_pipe_66_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	19 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_66_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_66_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_66_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_73_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_73_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_73_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_82_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_82_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_82_Sample/rr
      -- 
    ca_223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_66_inst_ack_1, ack => convTranspose_CP_39_elements(15)); -- 
    rr_259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(15), ack => RPIPE_ConvTranspose_input_pipe_82_inst_req_0); -- 
    rr_245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(15), ack => type_cast_73_inst_req_0); -- 
    -- CP-element group 16:  join  transition  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	11 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_68_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_68_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_68_Sample/req
      -- 
    req_231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(16), ack => WPIPE_ConvTranspose_output_pipe_68_inst_req_0); -- 
    convTranspose_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(11) & convTranspose_CP_39_elements(15);
      gj_convTranspose_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_68_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_68_update_start_
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_68_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_68_Sample/ack
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_68_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_68_Update/req
      -- 
    ack_232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_68_inst_ack_0, ack => convTranspose_CP_39_elements(17)); -- 
    req_236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(17), ack => WPIPE_ConvTranspose_output_pipe_68_inst_req_1); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	23 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_68_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_68_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_68_Update/ack
      -- 
    ack_237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_68_inst_ack_1, ack => convTranspose_CP_39_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_73_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_73_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_73_Sample/ra
      -- 
    ra_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_73_inst_ack_0, ack => convTranspose_CP_39_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	101 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_73_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_73_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_73_Update/ca
      -- 
    ca_251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_73_inst_ack_1, ack => convTranspose_CP_39_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_82_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_82_update_start_
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_82_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_82_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_82_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_82_Update/cr
      -- 
    ra_260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_82_inst_ack_0, ack => convTranspose_CP_39_elements(21)); -- 
    cr_264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(21), ack => RPIPE_ConvTranspose_input_pipe_82_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	28 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	26 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_82_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_82_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_82_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_89_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_89_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_89_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_97_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_97_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_97_Sample/rr
      -- 
    ca_265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_82_inst_ack_1, ack => convTranspose_CP_39_elements(22)); -- 
    rr_301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => RPIPE_ConvTranspose_input_pipe_97_inst_req_0); -- 
    rr_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => type_cast_89_inst_req_0); -- 
    -- CP-element group 23:  join  transition  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: 	18 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_84_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_84_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_84_Sample/req
      -- 
    req_273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(23), ack => WPIPE_ConvTranspose_output_pipe_84_inst_req_0); -- 
    convTranspose_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(22) & convTranspose_CP_39_elements(18);
      gj_convTranspose_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_84_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_84_update_start_
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_84_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_84_Sample/ack
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_84_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_84_Update/req
      -- 
    ack_274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_84_inst_ack_0, ack => convTranspose_CP_39_elements(24)); -- 
    req_278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(24), ack => WPIPE_ConvTranspose_output_pipe_84_inst_req_1); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	30 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_84_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_84_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_84_Update/ack
      -- 
    ack_279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_84_inst_ack_1, ack => convTranspose_CP_39_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	22 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_89_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_89_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_89_Sample/ra
      -- 
    ra_288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_89_inst_ack_0, ack => convTranspose_CP_39_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	101 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_89_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_89_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_89_Update/ca
      -- 
    ca_293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_89_inst_ack_1, ack => convTranspose_CP_39_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	22 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_97_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_97_update_start_
      -- CP-element group 28: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_97_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_97_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_97_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_97_Update/cr
      -- 
    ra_302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_97_inst_ack_0, ack => convTranspose_CP_39_elements(28)); -- 
    cr_306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(28), ack => RPIPE_ConvTranspose_input_pipe_97_inst_req_1); -- 
    -- CP-element group 29:  fork  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	33 
    -- CP-element group 29: 	30 
    -- CP-element group 29: 	35 
    -- CP-element group 29:  members (9) 
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_97_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_97_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_97_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_104_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_104_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_104_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_113_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_113_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_113_Sample/rr
      -- 
    ca_307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_97_inst_ack_1, ack => convTranspose_CP_39_elements(29)); -- 
    rr_343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(29), ack => RPIPE_ConvTranspose_input_pipe_113_inst_req_0); -- 
    rr_329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(29), ack => type_cast_104_inst_req_0); -- 
    -- CP-element group 30:  join  transition  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	25 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_99_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_99_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_99_Sample/req
      -- 
    req_315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(30), ack => WPIPE_ConvTranspose_output_pipe_99_inst_req_0); -- 
    convTranspose_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(25) & convTranspose_CP_39_elements(29);
      gj_convTranspose_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_99_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_99_update_start_
      -- CP-element group 31: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_99_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_99_Sample/ack
      -- CP-element group 31: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_99_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_99_Update/req
      -- 
    ack_316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_99_inst_ack_0, ack => convTranspose_CP_39_elements(31)); -- 
    req_320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(31), ack => WPIPE_ConvTranspose_output_pipe_99_inst_req_1); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	37 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_99_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_99_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_99_Update/ack
      -- 
    ack_321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_99_inst_ack_1, ack => convTranspose_CP_39_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	29 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_104_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_104_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_104_Sample/ra
      -- 
    ra_330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_104_inst_ack_0, ack => convTranspose_CP_39_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	0 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	104 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_104_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_104_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_104_Update/ca
      -- 
    ca_335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_104_inst_ack_1, ack => convTranspose_CP_39_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	29 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (6) 
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_113_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_113_update_start_
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_113_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_113_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_113_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_113_Update/cr
      -- 
    ra_344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_113_inst_ack_0, ack => convTranspose_CP_39_elements(35)); -- 
    cr_348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(35), ack => RPIPE_ConvTranspose_input_pipe_113_inst_req_1); -- 
    -- CP-element group 36:  fork  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	42 
    -- CP-element group 36: 	40 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (9) 
      -- CP-element group 36: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_113_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_113_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_113_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_120_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_120_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_120_Sample/rr
      -- CP-element group 36: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_128_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_128_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_128_Sample/rr
      -- 
    ca_349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_113_inst_ack_1, ack => convTranspose_CP_39_elements(36)); -- 
    rr_371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(36), ack => type_cast_120_inst_req_0); -- 
    rr_385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(36), ack => RPIPE_ConvTranspose_input_pipe_128_inst_req_0); -- 
    -- CP-element group 37:  join  transition  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	32 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_115_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_115_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_115_sample_start_
      -- 
    req_357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(37), ack => WPIPE_ConvTranspose_output_pipe_115_inst_req_0); -- 
    convTranspose_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(32) & convTranspose_CP_39_elements(36);
      gj_convTranspose_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_115_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_115_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_115_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_115_Update/req
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_115_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_115_update_start_
      -- 
    ack_358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_115_inst_ack_0, ack => convTranspose_CP_39_elements(38)); -- 
    req_362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(38), ack => WPIPE_ConvTranspose_output_pipe_115_inst_req_1); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	44 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_115_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_115_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_115_Update/ack
      -- 
    ack_363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_115_inst_ack_1, ack => convTranspose_CP_39_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	36 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_120_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_120_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_120_Sample/ra
      -- 
    ra_372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_120_inst_ack_0, ack => convTranspose_CP_39_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	0 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	104 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_120_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_120_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_120_Update/ca
      -- 
    ca_377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_120_inst_ack_1, ack => convTranspose_CP_39_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	36 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_128_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_128_update_start_
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_128_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_128_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_128_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_128_Update/cr
      -- 
    ra_386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_128_inst_ack_0, ack => convTranspose_CP_39_elements(42)); -- 
    cr_390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(42), ack => RPIPE_ConvTranspose_input_pipe_128_inst_req_1); -- 
    -- CP-element group 43:  fork  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	47 
    -- CP-element group 43: 	49 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_128_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_128_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_128_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_135_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_135_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_135_Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_144_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_144_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_144_Sample/rr
      -- 
    ca_391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_128_inst_ack_1, ack => convTranspose_CP_39_elements(43)); -- 
    rr_427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(43), ack => RPIPE_ConvTranspose_input_pipe_144_inst_req_0); -- 
    rr_413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(43), ack => type_cast_135_inst_req_0); -- 
    -- CP-element group 44:  join  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	39 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_130_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_130_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_130_Sample/req
      -- 
    req_399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(44), ack => WPIPE_ConvTranspose_output_pipe_130_inst_req_0); -- 
    convTranspose_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(39) & convTranspose_CP_39_elements(43);
      gj_convTranspose_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_130_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_130_update_start_
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_130_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_130_Sample/ack
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_130_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_130_Update/req
      -- 
    ack_400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_130_inst_ack_0, ack => convTranspose_CP_39_elements(45)); -- 
    req_404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(45), ack => WPIPE_ConvTranspose_output_pipe_130_inst_req_1); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	51 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_130_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_130_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_130_Update/ack
      -- 
    ack_405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_130_inst_ack_1, ack => convTranspose_CP_39_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	43 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_135_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_135_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_135_Sample/ra
      -- 
    ra_414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_135_inst_ack_0, ack => convTranspose_CP_39_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	107 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_135_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_135_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_135_Update/ca
      -- 
    ca_419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_135_inst_ack_1, ack => convTranspose_CP_39_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	43 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_144_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_144_update_start_
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_144_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_144_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_144_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_144_Update/cr
      -- 
    ra_428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_144_inst_ack_0, ack => convTranspose_CP_39_elements(49)); -- 
    cr_432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(49), ack => RPIPE_ConvTranspose_input_pipe_144_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	54 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	56 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_144_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_144_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_144_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_151_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_151_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_151_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_159_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_159_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_159_Sample/rr
      -- 
    ca_433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_144_inst_ack_1, ack => convTranspose_CP_39_elements(50)); -- 
    rr_469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => RPIPE_ConvTranspose_input_pipe_159_inst_req_0); -- 
    rr_455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => type_cast_151_inst_req_0); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	46 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_146_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_146_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_146_Sample/req
      -- 
    req_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(51), ack => WPIPE_ConvTranspose_output_pipe_146_inst_req_0); -- 
    convTranspose_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(46) & convTranspose_CP_39_elements(50);
      gj_convTranspose_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (6) 
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_146_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_146_update_start_
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_146_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_146_Sample/ack
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_146_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_146_Update/req
      -- 
    ack_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_146_inst_ack_0, ack => convTranspose_CP_39_elements(52)); -- 
    req_446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(52), ack => WPIPE_ConvTranspose_output_pipe_146_inst_req_1); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	58 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_146_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_146_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_146_Update/ack
      -- 
    ack_447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_146_inst_ack_1, ack => convTranspose_CP_39_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	50 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_151_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_151_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_151_Sample/ra
      -- 
    ra_456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_151_inst_ack_0, ack => convTranspose_CP_39_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	0 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	107 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_151_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_151_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_151_Update/ca
      -- 
    ca_461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_151_inst_ack_1, ack => convTranspose_CP_39_elements(55)); -- 
    -- CP-element group 56:  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	50 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (6) 
      -- CP-element group 56: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_159_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_159_update_start_
      -- CP-element group 56: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_159_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_159_Sample/ra
      -- CP-element group 56: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_159_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_159_Update/cr
      -- 
    ra_470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_159_inst_ack_0, ack => convTranspose_CP_39_elements(56)); -- 
    cr_474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(56), ack => RPIPE_ConvTranspose_input_pipe_159_inst_req_1); -- 
    -- CP-element group 57:  fork  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	61 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_159_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_159_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_159_Update/ca
      -- CP-element group 57: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_166_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_166_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_166_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_175_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_175_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_175_Sample/rr
      -- 
    ca_475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_159_inst_ack_1, ack => convTranspose_CP_39_elements(57)); -- 
    rr_497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(57), ack => type_cast_166_inst_req_0); -- 
    rr_511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(57), ack => RPIPE_ConvTranspose_input_pipe_175_inst_req_0); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	53 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_161_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_161_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_161_Sample/req
      -- 
    req_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(58), ack => WPIPE_ConvTranspose_output_pipe_161_inst_req_0); -- 
    convTranspose_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(53) & convTranspose_CP_39_elements(57);
      gj_convTranspose_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_161_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_161_update_start_
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_161_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_161_Sample/ack
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_161_Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_161_Update/req
      -- 
    ack_484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_161_inst_ack_0, ack => convTranspose_CP_39_elements(59)); -- 
    req_488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(59), ack => WPIPE_ConvTranspose_output_pipe_161_inst_req_1); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	65 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_161_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_161_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_161_Update/ack
      -- 
    ack_489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_161_inst_ack_1, ack => convTranspose_CP_39_elements(60)); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	57 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_166_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_166_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_166_Sample/ra
      -- 
    ra_498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_166_inst_ack_0, ack => convTranspose_CP_39_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	0 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	110 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_166_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_166_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_166_Update/ca
      -- 
    ca_503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_166_inst_ack_1, ack => convTranspose_CP_39_elements(62)); -- 
    -- CP-element group 63:  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_175_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_175_update_start_
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_175_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_175_Sample/ra
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_175_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_175_Update/cr
      -- 
    ra_512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_175_inst_ack_0, ack => convTranspose_CP_39_elements(63)); -- 
    cr_516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(63), ack => RPIPE_ConvTranspose_input_pipe_175_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	68 
    -- CP-element group 64: 	70 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (9) 
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_175_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_175_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_175_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_182_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_182_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_182_Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_190_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_190_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_190_Sample/rr
      -- 
    ca_517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_175_inst_ack_1, ack => convTranspose_CP_39_elements(64)); -- 
    rr_553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(64), ack => RPIPE_ConvTranspose_input_pipe_190_inst_req_0); -- 
    rr_539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(64), ack => type_cast_182_inst_req_0); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	60 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_177_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_177_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_177_Sample/req
      -- 
    req_525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(65), ack => WPIPE_ConvTranspose_output_pipe_177_inst_req_0); -- 
    convTranspose_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(60) & convTranspose_CP_39_elements(64);
      gj_convTranspose_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_177_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_177_update_start_
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_177_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_177_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_177_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_177_Update/req
      -- 
    ack_526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_177_inst_ack_0, ack => convTranspose_CP_39_elements(66)); -- 
    req_530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(66), ack => WPIPE_ConvTranspose_output_pipe_177_inst_req_1); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	72 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_177_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_177_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_177_Update/ack
      -- 
    ack_531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_177_inst_ack_1, ack => convTranspose_CP_39_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	64 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_182_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_182_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_182_Sample/ra
      -- 
    ra_540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_182_inst_ack_0, ack => convTranspose_CP_39_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	0 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	110 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_182_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_182_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_182_Update/ca
      -- 
    ca_545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_182_inst_ack_1, ack => convTranspose_CP_39_elements(69)); -- 
    -- CP-element group 70:  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	64 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (6) 
      -- CP-element group 70: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_190_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_190_update_start_
      -- CP-element group 70: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_190_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_190_Sample/ra
      -- CP-element group 70: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_190_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_190_Update/cr
      -- 
    ra_554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_190_inst_ack_0, ack => convTranspose_CP_39_elements(70)); -- 
    cr_558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(70), ack => RPIPE_ConvTranspose_input_pipe_190_inst_req_1); -- 
    -- CP-element group 71:  fork  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71: 	75 
    -- CP-element group 71: 	77 
    -- CP-element group 71:  members (9) 
      -- CP-element group 71: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_190_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_190_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_190_Update/ca
      -- CP-element group 71: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_197_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_197_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_197_Sample/rr
      -- CP-element group 71: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_206_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_206_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_206_Sample/rr
      -- 
    ca_559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_190_inst_ack_1, ack => convTranspose_CP_39_elements(71)); -- 
    rr_581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(71), ack => type_cast_197_inst_req_0); -- 
    rr_595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(71), ack => RPIPE_ConvTranspose_input_pipe_206_inst_req_0); -- 
    -- CP-element group 72:  join  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: 	67 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_192_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_192_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_192_Sample/req
      -- 
    req_567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(72), ack => WPIPE_ConvTranspose_output_pipe_192_inst_req_0); -- 
    convTranspose_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(71) & convTranspose_CP_39_elements(67);
      gj_convTranspose_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_192_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_192_update_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_192_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_192_Sample/ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_192_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_192_Update/req
      -- 
    ack_568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_192_inst_ack_0, ack => convTranspose_CP_39_elements(73)); -- 
    req_572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(73), ack => WPIPE_ConvTranspose_output_pipe_192_inst_req_1); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	79 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_192_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_192_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_192_Update/ack
      -- 
    ack_573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_192_inst_ack_1, ack => convTranspose_CP_39_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	71 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_197_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_197_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_197_Sample/ra
      -- 
    ra_582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_197_inst_ack_0, ack => convTranspose_CP_39_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	0 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	113 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_197_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_197_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_197_Update/ca
      -- 
    ca_587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_197_inst_ack_1, ack => convTranspose_CP_39_elements(76)); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	71 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_206_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_206_update_start_
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_206_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_206_Sample/ra
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_206_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_206_Update/cr
      -- 
    ra_596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_206_inst_ack_0, ack => convTranspose_CP_39_elements(77)); -- 
    cr_600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(77), ack => RPIPE_ConvTranspose_input_pipe_206_inst_req_1); -- 
    -- CP-element group 78:  fork  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	84 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	82 
    -- CP-element group 78:  members (9) 
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_206_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_206_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_206_Update/ca
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_213_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_213_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_213_Sample/rr
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_221_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_221_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_221_Sample/rr
      -- 
    ca_601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_206_inst_ack_1, ack => convTranspose_CP_39_elements(78)); -- 
    rr_623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(78), ack => type_cast_213_inst_req_0); -- 
    rr_637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(78), ack => RPIPE_ConvTranspose_input_pipe_221_inst_req_0); -- 
    -- CP-element group 79:  join  transition  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	74 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_208_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_208_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_208_Sample/req
      -- 
    req_609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(79), ack => WPIPE_ConvTranspose_output_pipe_208_inst_req_0); -- 
    convTranspose_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(74) & convTranspose_CP_39_elements(78);
      gj_convTranspose_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (6) 
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_208_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_208_update_start_
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_208_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_208_Sample/ack
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_208_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_208_Update/req
      -- 
    ack_610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_208_inst_ack_0, ack => convTranspose_CP_39_elements(80)); -- 
    req_614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(80), ack => WPIPE_ConvTranspose_output_pipe_208_inst_req_1); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	86 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_208_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_208_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_208_Update/ack
      -- 
    ack_615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_208_inst_ack_1, ack => convTranspose_CP_39_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	78 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_213_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_213_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_213_Sample/ra
      -- 
    ra_624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_213_inst_ack_0, ack => convTranspose_CP_39_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	0 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	113 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_213_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_213_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_213_Update/ca
      -- 
    ca_629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_213_inst_ack_1, ack => convTranspose_CP_39_elements(83)); -- 
    -- CP-element group 84:  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	78 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (6) 
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_221_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_221_update_start_
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_221_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_221_Sample/ra
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_221_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_221_Update/cr
      -- 
    ra_638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_221_inst_ack_0, ack => convTranspose_CP_39_elements(84)); -- 
    cr_642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(84), ack => RPIPE_ConvTranspose_input_pipe_221_inst_req_1); -- 
    -- CP-element group 85:  fork  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85: 	89 
    -- CP-element group 85: 	91 
    -- CP-element group 85:  members (9) 
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_221_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_221_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_221_Update/ca
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_228_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_228_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_228_Sample/rr
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_237_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_237_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_237_Sample/rr
      -- 
    ca_643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_221_inst_ack_1, ack => convTranspose_CP_39_elements(85)); -- 
    rr_665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(85), ack => type_cast_228_inst_req_0); -- 
    rr_679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(85), ack => RPIPE_ConvTranspose_input_pipe_237_inst_req_0); -- 
    -- CP-element group 86:  join  transition  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: 	81 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_223_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_223_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_223_Sample/req
      -- 
    req_651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(86), ack => WPIPE_ConvTranspose_output_pipe_223_inst_req_0); -- 
    convTranspose_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(85) & convTranspose_CP_39_elements(81);
      gj_convTranspose_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_223_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_223_update_start_
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_223_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_223_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_223_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_223_Update/req
      -- 
    ack_652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_223_inst_ack_0, ack => convTranspose_CP_39_elements(87)); -- 
    req_656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(87), ack => WPIPE_ConvTranspose_output_pipe_223_inst_req_1); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	93 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_223_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_223_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_223_Update/ack
      -- 
    ack_657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_223_inst_ack_1, ack => convTranspose_CP_39_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	85 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_228_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_228_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_228_Sample/ra
      -- 
    ra_666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_228_inst_ack_0, ack => convTranspose_CP_39_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	0 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	116 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_228_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_228_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_228_Update/ca
      -- 
    ca_671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_228_inst_ack_1, ack => convTranspose_CP_39_elements(90)); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	85 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_237_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_237_update_start_
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_237_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_237_Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_237_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_237_Update/cr
      -- 
    ra_680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_237_inst_ack_0, ack => convTranspose_CP_39_elements(91)); -- 
    cr_684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(91), ack => RPIPE_ConvTranspose_input_pipe_237_inst_req_1); -- 
    -- CP-element group 92:  fork  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92: 	96 
    -- CP-element group 92: 	119 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_237_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_237_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_237_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_244_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_244_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_244_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_305_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_305_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_305_Sample/rr
      -- 
    ca_685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_237_inst_ack_1, ack => convTranspose_CP_39_elements(92)); -- 
    rr_707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(92), ack => type_cast_244_inst_req_0); -- 
    rr_819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(92), ack => RPIPE_ConvTranspose_input_pipe_305_inst_req_0); -- 
    -- CP-element group 93:  join  transition  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	88 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_239_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_239_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_239_Sample/req
      -- 
    req_693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(93), ack => WPIPE_ConvTranspose_output_pipe_239_inst_req_0); -- 
    convTranspose_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(88) & convTranspose_CP_39_elements(92);
      gj_convTranspose_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_239_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_239_update_start_
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_239_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_239_Sample/ack
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_239_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_239_Update/req
      -- 
    ack_694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_239_inst_ack_0, ack => convTranspose_CP_39_elements(94)); -- 
    req_698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(94), ack => WPIPE_ConvTranspose_output_pipe_239_inst_req_1); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	121 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_239_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_239_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_239_Update/ack
      -- 
    ack_699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_239_inst_ack_1, ack => convTranspose_CP_39_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	92 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_244_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_244_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_244_Sample/ra
      -- 
    ra_708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_244_inst_ack_0, ack => convTranspose_CP_39_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	116 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_244_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_244_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_244_Update/ca
      -- 
    ca_713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_244_inst_ack_1, ack => convTranspose_CP_39_elements(97)); -- 
    -- CP-element group 98:  join  transition  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	6 
    -- CP-element group 98: 	13 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_253_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_253_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_253_Sample/rr
      -- 
    rr_721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(98), ack => type_cast_253_inst_req_0); -- 
    convTranspose_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(6) & convTranspose_CP_39_elements(13);
      gj_convTranspose_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_253_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_253_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_253_Sample/ra
      -- 
    ra_722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_253_inst_ack_0, ack => convTranspose_CP_39_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	0 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	189 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_253_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_253_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_253_Update/ca
      -- 
    ca_727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_253_inst_ack_1, ack => convTranspose_CP_39_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	27 
    -- CP-element group 101: 	20 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_257_sample_start_
      -- CP-element group 101: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_257_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_257_Sample/rr
      -- 
    rr_735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(101), ack => type_cast_257_inst_req_0); -- 
    convTranspose_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(27) & convTranspose_CP_39_elements(20);
      gj_convTranspose_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_257_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_257_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_257_Sample/ra
      -- 
    ra_736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_257_inst_ack_0, ack => convTranspose_CP_39_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	0 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	189 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_257_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_257_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_257_Update/ca
      -- 
    ca_741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_257_inst_ack_1, ack => convTranspose_CP_39_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	34 
    -- CP-element group 104: 	41 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_261_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_261_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_261_sample_start_
      -- 
    rr_749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(104), ack => type_cast_261_inst_req_0); -- 
    convTranspose_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(34) & convTranspose_CP_39_elements(41);
      gj_convTranspose_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_261_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_261_Sample/ra
      -- CP-element group 105: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_261_sample_completed_
      -- 
    ra_750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_261_inst_ack_0, ack => convTranspose_CP_39_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	0 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	189 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_261_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_261_Update/ca
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_261_update_completed_
      -- 
    ca_755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_261_inst_ack_1, ack => convTranspose_CP_39_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	55 
    -- CP-element group 107: 	48 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_275_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_275_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_275_Sample/rr
      -- 
    rr_763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(107), ack => type_cast_275_inst_req_0); -- 
    convTranspose_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(55) & convTranspose_CP_39_elements(48);
      gj_convTranspose_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_275_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_275_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_275_Sample/ra
      -- 
    ra_764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_275_inst_ack_0, ack => convTranspose_CP_39_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	0 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	189 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_275_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_275_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_275_Update/ca
      -- 
    ca_769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_275_inst_ack_1, ack => convTranspose_CP_39_elements(109)); -- 
    -- CP-element group 110:  join  transition  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	69 
    -- CP-element group 110: 	62 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_279_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_279_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_279_Sample/rr
      -- 
    rr_777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(110), ack => type_cast_279_inst_req_0); -- 
    convTranspose_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(69) & convTranspose_CP_39_elements(62);
      gj_convTranspose_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_279_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_279_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_279_Sample/ra
      -- 
    ra_778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_279_inst_ack_0, ack => convTranspose_CP_39_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	0 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	189 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_279_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_279_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_279_Update/ca
      -- 
    ca_783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_279_inst_ack_1, ack => convTranspose_CP_39_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	76 
    -- CP-element group 113: 	83 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_283_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_283_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_283_Sample/rr
      -- 
    rr_791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(113), ack => type_cast_283_inst_req_0); -- 
    convTranspose_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(76) & convTranspose_CP_39_elements(83);
      gj_convTranspose_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_283_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_283_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_283_Sample/ra
      -- 
    ra_792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_283_inst_ack_0, ack => convTranspose_CP_39_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	0 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	189 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_283_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_283_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_283_Update/ca
      -- 
    ca_797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_283_inst_ack_1, ack => convTranspose_CP_39_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	90 
    -- CP-element group 116: 	97 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_287_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_287_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_287_Sample/rr
      -- 
    rr_805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(116), ack => type_cast_287_inst_req_0); -- 
    convTranspose_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(90) & convTranspose_CP_39_elements(97);
      gj_convTranspose_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_287_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_287_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_287_Sample/ra
      -- 
    ra_806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_287_inst_ack_0, ack => convTranspose_CP_39_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	0 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	189 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_287_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_287_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_287_Update/ca
      -- 
    ca_811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_287_inst_ack_1, ack => convTranspose_CP_39_elements(118)); -- 
    -- CP-element group 119:  transition  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	92 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (6) 
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_305_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_305_update_start_
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_305_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_305_Sample/ra
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_305_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_305_Update/cr
      -- 
    ra_820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_305_inst_ack_0, ack => convTranspose_CP_39_elements(119)); -- 
    cr_824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(119), ack => RPIPE_ConvTranspose_input_pipe_305_inst_req_1); -- 
    -- CP-element group 120:  fork  transition  input  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120: 	124 
    -- CP-element group 120: 	126 
    -- CP-element group 120:  members (9) 
      -- CP-element group 120: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_305_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_305_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_305_Update/ca
      -- CP-element group 120: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_312_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_312_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_312_Sample/rr
      -- CP-element group 120: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_321_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_321_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_321_Sample/rr
      -- 
    ca_825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_305_inst_ack_1, ack => convTranspose_CP_39_elements(120)); -- 
    rr_847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(120), ack => type_cast_312_inst_req_0); -- 
    rr_861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(120), ack => RPIPE_ConvTranspose_input_pipe_321_inst_req_0); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	95 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_307_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_307_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_307_Sample/req
      -- 
    req_833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(121), ack => WPIPE_ConvTranspose_output_pipe_307_inst_req_0); -- 
    convTranspose_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(95) & convTranspose_CP_39_elements(120);
      gj_convTranspose_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  transition  input  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (6) 
      -- CP-element group 122: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_307_sample_completed_
      -- CP-element group 122: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_307_update_start_
      -- CP-element group 122: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_307_Sample/$exit
      -- CP-element group 122: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_307_Sample/ack
      -- CP-element group 122: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_307_Update/$entry
      -- CP-element group 122: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_307_Update/req
      -- 
    ack_834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_307_inst_ack_0, ack => convTranspose_CP_39_elements(122)); -- 
    req_838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(122), ack => WPIPE_ConvTranspose_output_pipe_307_inst_req_1); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	128 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_307_update_completed_
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_307_Update/$exit
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_307_Update/ack
      -- 
    ack_839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_307_inst_ack_1, ack => convTranspose_CP_39_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	120 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_312_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_312_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_312_Sample/ra
      -- 
    ra_848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_312_inst_ack_0, ack => convTranspose_CP_39_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	0 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	189 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_312_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_312_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_312_Update/ca
      -- 
    ca_853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_312_inst_ack_1, ack => convTranspose_CP_39_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	120 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (6) 
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_321_sample_completed_
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_321_update_start_
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_321_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_321_Sample/ra
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_321_Update/$entry
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_321_Update/cr
      -- 
    ra_862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_321_inst_ack_0, ack => convTranspose_CP_39_elements(126)); -- 
    cr_866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(126), ack => RPIPE_ConvTranspose_input_pipe_321_inst_req_1); -- 
    -- CP-element group 127:  fork  transition  input  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	131 
    -- CP-element group 127: 	133 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (9) 
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_321_update_completed_
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_321_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_321_Update/ca
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_328_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_328_Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_328_Sample/rr
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_336_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_336_Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_336_Sample/rr
      -- 
    ca_867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_321_inst_ack_1, ack => convTranspose_CP_39_elements(127)); -- 
    rr_889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(127), ack => type_cast_328_inst_req_0); -- 
    rr_903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(127), ack => RPIPE_ConvTranspose_input_pipe_336_inst_req_0); -- 
    -- CP-element group 128:  join  transition  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	123 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_323_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_323_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_323_Sample/req
      -- 
    req_875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(128), ack => WPIPE_ConvTranspose_output_pipe_323_inst_req_0); -- 
    convTranspose_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(123) & convTranspose_CP_39_elements(127);
      gj_convTranspose_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_323_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_323_update_start_
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_323_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_323_Sample/ack
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_323_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_323_Update/req
      -- 
    ack_876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_323_inst_ack_0, ack => convTranspose_CP_39_elements(129)); -- 
    req_880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(129), ack => WPIPE_ConvTranspose_output_pipe_323_inst_req_1); -- 
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	135 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_323_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_323_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_323_Update/ack
      -- 
    ack_881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_323_inst_ack_1, ack => convTranspose_CP_39_elements(130)); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	127 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_328_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_328_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_328_Sample/ra
      -- 
    ra_890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_328_inst_ack_0, ack => convTranspose_CP_39_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	0 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	189 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_328_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_328_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_328_Update/ca
      -- 
    ca_895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_328_inst_ack_1, ack => convTranspose_CP_39_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	127 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_336_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_336_update_start_
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_336_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_336_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_336_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_336_Update/cr
      -- 
    ra_904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_336_inst_ack_0, ack => convTranspose_CP_39_elements(133)); -- 
    cr_908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(133), ack => RPIPE_ConvTranspose_input_pipe_336_inst_req_1); -- 
    -- CP-element group 134:  fork  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	138 
    -- CP-element group 134: 	140 
    -- CP-element group 134: 	135 
    -- CP-element group 134:  members (9) 
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_352_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_336_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_336_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_336_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_343_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_343_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_343_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_352_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_352_Sample/$entry
      -- 
    ca_909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_336_inst_ack_1, ack => convTranspose_CP_39_elements(134)); -- 
    rr_931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(134), ack => type_cast_343_inst_req_0); -- 
    rr_945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(134), ack => RPIPE_ConvTranspose_input_pipe_352_inst_req_0); -- 
    -- CP-element group 135:  join  transition  output  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	130 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_338_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_338_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_338_Sample/req
      -- 
    req_917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(135), ack => WPIPE_ConvTranspose_output_pipe_338_inst_req_0); -- 
    convTranspose_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(130) & convTranspose_CP_39_elements(134);
      gj_convTranspose_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  transition  input  output  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (6) 
      -- CP-element group 136: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_338_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_338_update_start_
      -- CP-element group 136: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_338_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_338_Sample/ack
      -- CP-element group 136: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_338_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_338_Update/req
      -- 
    ack_918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_338_inst_ack_0, ack => convTranspose_CP_39_elements(136)); -- 
    req_922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(136), ack => WPIPE_ConvTranspose_output_pipe_338_inst_req_1); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	142 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_338_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_338_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_338_Update/ack
      -- 
    ack_923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_338_inst_ack_1, ack => convTranspose_CP_39_elements(137)); -- 
    -- CP-element group 138:  transition  input  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	134 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_343_sample_completed_
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_343_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_343_Sample/ra
      -- 
    ra_932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_343_inst_ack_0, ack => convTranspose_CP_39_elements(138)); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	0 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	189 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_343_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_343_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_343_Update/ca
      -- 
    ca_937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_343_inst_ack_1, ack => convTranspose_CP_39_elements(139)); -- 
    -- CP-element group 140:  transition  input  output  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	134 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	141 
    -- CP-element group 140:  members (6) 
      -- CP-element group 140: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_352_Update/$entry
      -- CP-element group 140: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_352_Update/cr
      -- CP-element group 140: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_352_Sample/ra
      -- CP-element group 140: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_352_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_352_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_352_update_start_
      -- 
    ra_946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_352_inst_ack_0, ack => convTranspose_CP_39_elements(140)); -- 
    cr_950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(140), ack => RPIPE_ConvTranspose_input_pipe_352_inst_req_1); -- 
    -- CP-element group 141:  fork  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	140 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	145 
    -- CP-element group 141: 	147 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (9) 
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_352_Update/ca
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_352_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_367_Sample/rr
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_367_Sample/$entry
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_367_sample_start_
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_359_Sample/rr
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_359_Sample/$entry
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_359_sample_start_
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_352_update_completed_
      -- 
    ca_951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_352_inst_ack_1, ack => convTranspose_CP_39_elements(141)); -- 
    rr_987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(141), ack => RPIPE_ConvTranspose_input_pipe_367_inst_req_0); -- 
    rr_973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(141), ack => type_cast_359_inst_req_0); -- 
    -- CP-element group 142:  join  transition  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	137 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_354_Sample/req
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_354_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_354_sample_start_
      -- 
    req_959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(142), ack => WPIPE_ConvTranspose_output_pipe_354_inst_req_0); -- 
    convTranspose_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(137) & convTranspose_CP_39_elements(141);
      gj_convTranspose_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143:  members (6) 
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_354_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_354_update_start_
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_354_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_354_Update/req
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_354_Update/$entry
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_354_Sample/ack
      -- 
    ack_960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_354_inst_ack_0, ack => convTranspose_CP_39_elements(143)); -- 
    req_964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(143), ack => WPIPE_ConvTranspose_output_pipe_354_inst_req_1); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	149 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_354_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_354_Update/ack
      -- CP-element group 144: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_354_Update/$exit
      -- 
    ack_965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_354_inst_ack_1, ack => convTranspose_CP_39_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	141 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_359_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_359_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_359_sample_completed_
      -- 
    ra_974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_359_inst_ack_0, ack => convTranspose_CP_39_elements(145)); -- 
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	0 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	189 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_359_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_359_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_359_update_completed_
      -- 
    ca_979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_359_inst_ack_1, ack => convTranspose_CP_39_elements(146)); -- 
    -- CP-element group 147:  transition  input  output  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	141 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	148 
    -- CP-element group 147:  members (6) 
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_367_Update/cr
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_367_Update/$entry
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_367_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_367_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_367_update_start_
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_367_sample_completed_
      -- 
    ra_988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_367_inst_ack_0, ack => convTranspose_CP_39_elements(147)); -- 
    cr_992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(147), ack => RPIPE_ConvTranspose_input_pipe_367_inst_req_1); -- 
    -- CP-element group 148:  fork  transition  input  output  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	147 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	154 
    -- CP-element group 148: 	149 
    -- CP-element group 148: 	152 
    -- CP-element group 148:  members (9) 
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_383_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_383_Sample/rr
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_383_Sample/$entry
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_374_Sample/rr
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_374_Sample/$entry
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_374_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_367_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_367_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_367_update_completed_
      -- 
    ca_993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_367_inst_ack_1, ack => convTranspose_CP_39_elements(148)); -- 
    rr_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(148), ack => RPIPE_ConvTranspose_input_pipe_383_inst_req_0); -- 
    rr_1015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(148), ack => type_cast_374_inst_req_0); -- 
    -- CP-element group 149:  join  transition  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	148 
    -- CP-element group 149: 	144 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_369_Sample/req
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_369_Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_369_sample_start_
      -- 
    req_1001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(149), ack => WPIPE_ConvTranspose_output_pipe_369_inst_req_0); -- 
    convTranspose_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(148) & convTranspose_CP_39_elements(144);
      gj_convTranspose_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150:  members (6) 
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_369_Update/req
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_369_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_369_Sample/ack
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_369_Sample/$exit
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_369_update_start_
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_369_sample_completed_
      -- 
    ack_1002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_369_inst_ack_0, ack => convTranspose_CP_39_elements(150)); -- 
    req_1006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(150), ack => WPIPE_ConvTranspose_output_pipe_369_inst_req_1); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	156 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_369_Update/ack
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_369_Update/$exit
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_369_update_completed_
      -- 
    ack_1007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_369_inst_ack_1, ack => convTranspose_CP_39_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	148 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_374_Sample/ra
      -- CP-element group 152: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_374_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_374_sample_completed_
      -- 
    ra_1016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_374_inst_ack_0, ack => convTranspose_CP_39_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	0 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	189 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_374_Update/ca
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_374_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_374_update_completed_
      -- 
    ca_1021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_374_inst_ack_1, ack => convTranspose_CP_39_elements(153)); -- 
    -- CP-element group 154:  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	148 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (6) 
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_383_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_383_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_383_Sample/ra
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_383_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_383_update_start_
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_383_sample_completed_
      -- 
    ra_1030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_383_inst_ack_0, ack => convTranspose_CP_39_elements(154)); -- 
    cr_1034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(154), ack => RPIPE_ConvTranspose_input_pipe_383_inst_req_1); -- 
    -- CP-element group 155:  fork  transition  input  output  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: 	159 
    -- CP-element group 155: 	161 
    -- CP-element group 155:  members (9) 
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_390_Sample/rr
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_383_Update/ca
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_383_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_383_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_390_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_390_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_398_Sample/rr
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_398_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_398_sample_start_
      -- 
    ca_1035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_383_inst_ack_1, ack => convTranspose_CP_39_elements(155)); -- 
    rr_1057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(155), ack => type_cast_390_inst_req_0); -- 
    rr_1071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(155), ack => RPIPE_ConvTranspose_input_pipe_398_inst_req_0); -- 
    -- CP-element group 156:  join  transition  output  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: 	151 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	157 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_385_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_385_Sample/req
      -- CP-element group 156: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_385_Sample/$entry
      -- 
    req_1043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(156), ack => WPIPE_ConvTranspose_output_pipe_385_inst_req_0); -- 
    convTranspose_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(155) & convTranspose_CP_39_elements(151);
      gj_convTranspose_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	156 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_385_update_start_
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_385_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_385_Update/req
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_385_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_385_Sample/ack
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_385_Sample/$exit
      -- 
    ack_1044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_385_inst_ack_0, ack => convTranspose_CP_39_elements(157)); -- 
    req_1048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(157), ack => WPIPE_ConvTranspose_output_pipe_385_inst_req_1); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	163 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_385_Update/ack
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_385_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_385_update_completed_
      -- 
    ack_1049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_385_inst_ack_1, ack => convTranspose_CP_39_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	155 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_390_Sample/ra
      -- CP-element group 159: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_390_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_390_Sample/$exit
      -- 
    ra_1058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_390_inst_ack_0, ack => convTranspose_CP_39_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	0 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	189 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_390_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_390_Update/ca
      -- CP-element group 160: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_390_Update/$exit
      -- 
    ca_1063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_390_inst_ack_1, ack => convTranspose_CP_39_elements(160)); -- 
    -- CP-element group 161:  transition  input  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	155 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (6) 
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_398_update_start_
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_398_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_398_Update/cr
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_398_Update/$entry
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_398_Sample/ra
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_398_Sample/$exit
      -- 
    ra_1072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_398_inst_ack_0, ack => convTranspose_CP_39_elements(161)); -- 
    cr_1076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(161), ack => RPIPE_ConvTranspose_input_pipe_398_inst_req_1); -- 
    -- CP-element group 162:  fork  transition  input  output  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162: 	166 
    -- CP-element group 162: 	168 
    -- CP-element group 162:  members (9) 
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_405_Sample/rr
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_405_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_405_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_414_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_398_Update/ca
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_398_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_414_Sample/rr
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_398_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_414_sample_start_
      -- 
    ca_1077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_398_inst_ack_1, ack => convTranspose_CP_39_elements(162)); -- 
    rr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(162), ack => type_cast_405_inst_req_0); -- 
    rr_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(162), ack => RPIPE_ConvTranspose_input_pipe_414_inst_req_0); -- 
    -- CP-element group 163:  join  transition  output  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	158 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_400_Sample/req
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_400_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_400_sample_start_
      -- 
    req_1085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(163), ack => WPIPE_ConvTranspose_output_pipe_400_inst_req_0); -- 
    convTranspose_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(158) & convTranspose_CP_39_elements(162);
      gj_convTranspose_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  transition  input  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164:  members (6) 
      -- CP-element group 164: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_400_Update/req
      -- CP-element group 164: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_400_Update/$entry
      -- CP-element group 164: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_400_Sample/ack
      -- CP-element group 164: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_400_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_400_update_start_
      -- CP-element group 164: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_400_sample_completed_
      -- 
    ack_1086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_400_inst_ack_0, ack => convTranspose_CP_39_elements(164)); -- 
    req_1090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(164), ack => WPIPE_ConvTranspose_output_pipe_400_inst_req_1); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	170 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_400_Update/ack
      -- CP-element group 165: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_400_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_400_update_completed_
      -- 
    ack_1091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_400_inst_ack_1, ack => convTranspose_CP_39_elements(165)); -- 
    -- CP-element group 166:  transition  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	162 
    -- CP-element group 166: successors 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_405_Sample/ra
      -- CP-element group 166: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_405_Sample/$exit
      -- CP-element group 166: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_405_sample_completed_
      -- 
    ra_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_405_inst_ack_0, ack => convTranspose_CP_39_elements(166)); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	0 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	189 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_405_Update/ca
      -- CP-element group 167: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_405_Update/$exit
      -- CP-element group 167: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_405_update_completed_
      -- 
    ca_1105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_405_inst_ack_1, ack => convTranspose_CP_39_elements(167)); -- 
    -- CP-element group 168:  transition  input  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	162 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (6) 
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_414_update_start_
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_414_Update/cr
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_414_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_414_Sample/ra
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_414_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_414_sample_completed_
      -- 
    ra_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_414_inst_ack_0, ack => convTranspose_CP_39_elements(168)); -- 
    cr_1118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(168), ack => RPIPE_ConvTranspose_input_pipe_414_inst_req_1); -- 
    -- CP-element group 169:  fork  transition  input  output  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169: 	173 
    -- CP-element group 169: 	175 
    -- CP-element group 169:  members (9) 
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_421_sample_start_
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_414_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_429_Sample/rr
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_429_Sample/$entry
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_429_sample_start_
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_414_Update/ca
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_414_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_421_Sample/rr
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_421_Sample/$entry
      -- 
    ca_1119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_414_inst_ack_1, ack => convTranspose_CP_39_elements(169)); -- 
    rr_1141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(169), ack => type_cast_421_inst_req_0); -- 
    rr_1155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(169), ack => RPIPE_ConvTranspose_input_pipe_429_inst_req_0); -- 
    -- CP-element group 170:  join  transition  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	165 
    -- CP-element group 170: 	169 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_416_Sample/req
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_416_Sample/$entry
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_416_sample_start_
      -- 
    req_1127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(170), ack => WPIPE_ConvTranspose_output_pipe_416_inst_req_0); -- 
    convTranspose_cp_element_group_170: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_170"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(165) & convTranspose_CP_39_elements(169);
      gj_convTranspose_cp_element_group_170 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(170), clk => clk, reset => reset); --
    end block;
    -- CP-element group 171:  transition  input  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171:  members (6) 
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_416_Update/req
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_416_Update/$entry
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_416_Sample/ack
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_416_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_416_update_start_
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_416_sample_completed_
      -- 
    ack_1128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_416_inst_ack_0, ack => convTranspose_CP_39_elements(171)); -- 
    req_1132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(171), ack => WPIPE_ConvTranspose_output_pipe_416_inst_req_1); -- 
    -- CP-element group 172:  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	177 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_416_Update/ack
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_416_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_416_update_completed_
      -- 
    ack_1133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_416_inst_ack_1, ack => convTranspose_CP_39_elements(172)); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	169 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_421_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_421_Sample/ra
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_421_Sample/$exit
      -- 
    ra_1142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_421_inst_ack_0, ack => convTranspose_CP_39_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	0 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	189 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_421_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_421_Update/ca
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_421_Update/$exit
      -- 
    ca_1147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_421_inst_ack_1, ack => convTranspose_CP_39_elements(174)); -- 
    -- CP-element group 175:  transition  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	169 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (6) 
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_429_Update/cr
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_429_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_429_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_429_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_429_update_start_
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_429_sample_completed_
      -- 
    ra_1156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_429_inst_ack_0, ack => convTranspose_CP_39_elements(175)); -- 
    cr_1160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(175), ack => RPIPE_ConvTranspose_input_pipe_429_inst_req_1); -- 
    -- CP-element group 176:  fork  transition  input  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176: 	180 
    -- CP-element group 176: 	182 
    -- CP-element group 176:  members (9) 
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_436_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_445_Sample/rr
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_429_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_429_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_445_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_429_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_445_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_436_Sample/rr
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_436_Sample/$entry
      -- 
    ca_1161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_429_inst_ack_1, ack => convTranspose_CP_39_elements(176)); -- 
    rr_1183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(176), ack => type_cast_436_inst_req_0); -- 
    rr_1197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(176), ack => RPIPE_ConvTranspose_input_pipe_445_inst_req_0); -- 
    -- CP-element group 177:  join  transition  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	172 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_431_Sample/req
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_431_Sample/$entry
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_431_sample_start_
      -- 
    req_1169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(177), ack => WPIPE_ConvTranspose_output_pipe_431_inst_req_0); -- 
    convTranspose_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(172) & convTranspose_CP_39_elements(176);
      gj_convTranspose_cp_element_group_177 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (6) 
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_431_Update/req
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_431_Update/$entry
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_431_Sample/ack
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_431_Sample/$exit
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_431_update_start_
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_431_sample_completed_
      -- 
    ack_1170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_431_inst_ack_0, ack => convTranspose_CP_39_elements(178)); -- 
    req_1174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(178), ack => WPIPE_ConvTranspose_output_pipe_431_inst_req_1); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	184 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_431_Update/ack
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_431_Update/$exit
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_431_update_completed_
      -- 
    ack_1175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_431_inst_ack_1, ack => convTranspose_CP_39_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	176 
    -- CP-element group 180: successors 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_436_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_436_Sample/ra
      -- CP-element group 180: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_436_Sample/$exit
      -- 
    ra_1184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_436_inst_ack_0, ack => convTranspose_CP_39_elements(180)); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	0 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	189 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_436_Update/ca
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_436_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_436_update_completed_
      -- 
    ca_1189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_436_inst_ack_1, ack => convTranspose_CP_39_elements(181)); -- 
    -- CP-element group 182:  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	176 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182:  members (6) 
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_445_Update/cr
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_445_Update/$entry
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_445_Sample/ra
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_445_Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_445_update_start_
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_445_sample_completed_
      -- 
    ra_1198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_445_inst_ack_0, ack => convTranspose_CP_39_elements(182)); -- 
    cr_1202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(182), ack => RPIPE_ConvTranspose_input_pipe_445_inst_req_1); -- 
    -- CP-element group 183:  fork  transition  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183: 	187 
    -- CP-element group 183:  members (6) 
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_452_sample_start_
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_452_Sample/rr
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_452_Sample/$entry
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_445_Update/ca
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_445_Update/$exit
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/RPIPE_ConvTranspose_input_pipe_445_update_completed_
      -- 
    ca_1203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_445_inst_ack_1, ack => convTranspose_CP_39_elements(183)); -- 
    rr_1225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(183), ack => type_cast_452_inst_req_0); -- 
    -- CP-element group 184:  join  transition  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	179 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_447_Sample/req
      -- CP-element group 184: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_447_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_447_sample_start_
      -- 
    req_1211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(184), ack => WPIPE_ConvTranspose_output_pipe_447_inst_req_0); -- 
    convTranspose_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(179) & convTranspose_CP_39_elements(183);
      gj_convTranspose_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  transition  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (6) 
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_447_Update/req
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_447_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_447_Sample/ack
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_447_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_447_update_start_
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_447_sample_completed_
      -- 
    ack_1212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_447_inst_ack_0, ack => convTranspose_CP_39_elements(185)); -- 
    req_1216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(185), ack => WPIPE_ConvTranspose_output_pipe_447_inst_req_1); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	189 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_447_Update/ack
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_447_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/WPIPE_ConvTranspose_output_pipe_447_update_completed_
      -- 
    ack_1217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_447_inst_ack_1, ack => convTranspose_CP_39_elements(186)); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	183 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_452_Sample/ra
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_452_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_452_sample_completed_
      -- 
    ra_1226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_452_inst_ack_0, ack => convTranspose_CP_39_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	0 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_452_Update/ca
      -- CP-element group 188: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_452_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/type_cast_452_update_completed_
      -- 
    ca_1231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_452_inst_ack_1, ack => convTranspose_CP_39_elements(188)); -- 
    -- CP-element group 189:  branch  join  transition  place  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	153 
    -- CP-element group 189: 	160 
    -- CP-element group 189: 	167 
    -- CP-element group 189: 	174 
    -- CP-element group 189: 	181 
    -- CP-element group 189: 	186 
    -- CP-element group 189: 	188 
    -- CP-element group 189: 	100 
    -- CP-element group 189: 	146 
    -- CP-element group 189: 	139 
    -- CP-element group 189: 	112 
    -- CP-element group 189: 	115 
    -- CP-element group 189: 	118 
    -- CP-element group 189: 	103 
    -- CP-element group 189: 	106 
    -- CP-element group 189: 	109 
    -- CP-element group 189: 	132 
    -- CP-element group 189: 	125 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (10) 
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465__exit__
      -- CP-element group 189: 	 branch_block_stmt_33/if_stmt_466__entry__
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_465/$exit
      -- CP-element group 189: 	 branch_block_stmt_33/if_stmt_466_else_link/$entry
      -- CP-element group 189: 	 branch_block_stmt_33/if_stmt_466_if_link/$entry
      -- CP-element group 189: 	 branch_block_stmt_33/R_cmp575_467_place
      -- CP-element group 189: 	 branch_block_stmt_33/if_stmt_466_eval_test/branch_req
      -- CP-element group 189: 	 branch_block_stmt_33/if_stmt_466_eval_test/$exit
      -- CP-element group 189: 	 branch_block_stmt_33/if_stmt_466_eval_test/$entry
      -- CP-element group 189: 	 branch_block_stmt_33/if_stmt_466_dead_link/$entry
      -- 
    branch_req_1239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(189), ack => if_stmt_466_branch_req_0); -- 
    convTranspose_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 17) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1);
      constant place_markings: IntegerArray(0 to 17)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0);
      constant place_delays: IntegerArray(0 to 17) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 18); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(153) & convTranspose_CP_39_elements(160) & convTranspose_CP_39_elements(167) & convTranspose_CP_39_elements(174) & convTranspose_CP_39_elements(181) & convTranspose_CP_39_elements(186) & convTranspose_CP_39_elements(188) & convTranspose_CP_39_elements(100) & convTranspose_CP_39_elements(146) & convTranspose_CP_39_elements(139) & convTranspose_CP_39_elements(112) & convTranspose_CP_39_elements(115) & convTranspose_CP_39_elements(118) & convTranspose_CP_39_elements(103) & convTranspose_CP_39_elements(106) & convTranspose_CP_39_elements(109) & convTranspose_CP_39_elements(132) & convTranspose_CP_39_elements(125);
      gj_convTranspose_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 18, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	194 
    -- CP-element group 190: 	195 
    -- CP-element group 190:  members (18) 
      -- CP-element group 190: 	 branch_block_stmt_33/merge_stmt_487__exit__
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_493_to_assign_stmt_522__entry__
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_493_to_assign_stmt_522/type_cast_508_Update/cr
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_493_to_assign_stmt_522/type_cast_508_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_493_to_assign_stmt_522/type_cast_508_Sample/rr
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_493_to_assign_stmt_522/type_cast_508_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_493_to_assign_stmt_522/type_cast_508_update_start_
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_493_to_assign_stmt_522/type_cast_508_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_493_to_assign_stmt_522/$entry
      -- CP-element group 190: 	 branch_block_stmt_33/entry_bbx_xnph577
      -- CP-element group 190: 	 branch_block_stmt_33/if_stmt_466_if_link/if_choice_transition
      -- CP-element group 190: 	 branch_block_stmt_33/if_stmt_466_if_link/$exit
      -- CP-element group 190: 	 branch_block_stmt_33/entry_bbx_xnph577_PhiReq/$entry
      -- CP-element group 190: 	 branch_block_stmt_33/entry_bbx_xnph577_PhiReq/$exit
      -- CP-element group 190: 	 branch_block_stmt_33/merge_stmt_487_PhiReqMerge
      -- CP-element group 190: 	 branch_block_stmt_33/merge_stmt_487_PhiAck/$entry
      -- CP-element group 190: 	 branch_block_stmt_33/merge_stmt_487_PhiAck/$exit
      -- CP-element group 190: 	 branch_block_stmt_33/merge_stmt_487_PhiAck/dummy
      -- 
    if_choice_transition_1244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_466_branch_ack_1, ack => convTranspose_CP_39_elements(190)); -- 
    cr_1288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(190), ack => type_cast_508_inst_req_1); -- 
    rr_1283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(190), ack => type_cast_508_inst_req_0); -- 
    -- CP-element group 191:  transition  place  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	515 
    -- CP-element group 191:  members (5) 
      -- CP-element group 191: 	 branch_block_stmt_33/entry_forx_xcond302x_xpreheader
      -- CP-element group 191: 	 branch_block_stmt_33/if_stmt_466_else_link/else_choice_transition
      -- CP-element group 191: 	 branch_block_stmt_33/if_stmt_466_else_link/$exit
      -- CP-element group 191: 	 branch_block_stmt_33/entry_forx_xcond302x_xpreheader_PhiReq/$entry
      -- CP-element group 191: 	 branch_block_stmt_33/entry_forx_xcond302x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_1248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_466_branch_ack_0, ack => convTranspose_CP_39_elements(191)); -- 
    -- CP-element group 192:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	515 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	261 
    -- CP-element group 192: 	262 
    -- CP-element group 192:  members (18) 
      -- CP-element group 192: 	 branch_block_stmt_33/merge_stmt_718__exit__
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_724_to_assign_stmt_753__entry__
      -- CP-element group 192: 	 branch_block_stmt_33/if_stmt_481_if_link/if_choice_transition
      -- CP-element group 192: 	 branch_block_stmt_33/forx_xcond302x_xpreheader_bbx_xnph573
      -- CP-element group 192: 	 branch_block_stmt_33/if_stmt_481_if_link/$exit
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_724_to_assign_stmt_753/$entry
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_724_to_assign_stmt_753/type_cast_739_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_724_to_assign_stmt_753/type_cast_739_update_start_
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_724_to_assign_stmt_753/type_cast_739_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_724_to_assign_stmt_753/type_cast_739_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_724_to_assign_stmt_753/type_cast_739_Update/$entry
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_724_to_assign_stmt_753/type_cast_739_Update/cr
      -- CP-element group 192: 	 branch_block_stmt_33/forx_xcond302x_xpreheader_bbx_xnph573_PhiReq/$entry
      -- CP-element group 192: 	 branch_block_stmt_33/forx_xcond302x_xpreheader_bbx_xnph573_PhiReq/$exit
      -- CP-element group 192: 	 branch_block_stmt_33/merge_stmt_718_PhiReqMerge
      -- CP-element group 192: 	 branch_block_stmt_33/merge_stmt_718_PhiAck/$entry
      -- CP-element group 192: 	 branch_block_stmt_33/merge_stmt_718_PhiAck/$exit
      -- CP-element group 192: 	 branch_block_stmt_33/merge_stmt_718_PhiAck/dummy
      -- 
    if_choice_transition_1266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_481_branch_ack_1, ack => convTranspose_CP_39_elements(192)); -- 
    rr_1754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(192), ack => type_cast_739_inst_req_0); -- 
    cr_1759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(192), ack => type_cast_739_inst_req_1); -- 
    -- CP-element group 193:  transition  place  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	515 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	528 
    -- CP-element group 193:  members (5) 
      -- CP-element group 193: 	 branch_block_stmt_33/if_stmt_481_else_link/$exit
      -- CP-element group 193: 	 branch_block_stmt_33/forx_xcond302x_xpreheader_forx_xend394
      -- CP-element group 193: 	 branch_block_stmt_33/if_stmt_481_else_link/else_choice_transition
      -- CP-element group 193: 	 branch_block_stmt_33/forx_xcond302x_xpreheader_forx_xend394_PhiReq/$entry
      -- CP-element group 193: 	 branch_block_stmt_33/forx_xcond302x_xpreheader_forx_xend394_PhiReq/$exit
      -- 
    else_choice_transition_1270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_481_branch_ack_0, ack => convTranspose_CP_39_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	190 
    -- CP-element group 194: successors 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_493_to_assign_stmt_522/type_cast_508_Sample/ra
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_493_to_assign_stmt_522/type_cast_508_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_493_to_assign_stmt_522/type_cast_508_sample_completed_
      -- 
    ra_1284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_508_inst_ack_0, ack => convTranspose_CP_39_elements(194)); -- 
    -- CP-element group 195:  transition  place  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	190 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	516 
    -- CP-element group 195:  members (9) 
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_493_to_assign_stmt_522__exit__
      -- CP-element group 195: 	 branch_block_stmt_33/bbx_xnph577_forx_xbody
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_493_to_assign_stmt_522/type_cast_508_Update/ca
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_493_to_assign_stmt_522/type_cast_508_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_493_to_assign_stmt_522/type_cast_508_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_493_to_assign_stmt_522/$exit
      -- CP-element group 195: 	 branch_block_stmt_33/bbx_xnph577_forx_xbody_PhiReq/$entry
      -- CP-element group 195: 	 branch_block_stmt_33/bbx_xnph577_forx_xbody_PhiReq/phi_stmt_525/$entry
      -- CP-element group 195: 	 branch_block_stmt_33/bbx_xnph577_forx_xbody_PhiReq/phi_stmt_525/phi_stmt_525_sources/$entry
      -- 
    ca_1289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_508_inst_ack_1, ack => convTranspose_CP_39_elements(195)); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	521 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	258 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_final_index_sum_regn_sample_complete
      -- CP-element group 196: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_final_index_sum_regn_Sample/ack
      -- CP-element group 196: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_final_index_sum_regn_Sample/$exit
      -- 
    ack_1318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_537_index_offset_ack_0, ack => convTranspose_CP_39_elements(196)); -- 
    -- CP-element group 197:  transition  input  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	521 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (11) 
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/addr_of_538_request/req
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/addr_of_538_request/$entry
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_base_plus_offset/$exit
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_base_plus_offset/sum_rename_ack
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_base_plus_offset/sum_rename_req
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/addr_of_538_sample_start_
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_base_plus_offset/$entry
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_final_index_sum_regn_Update/ack
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_offset_calculated
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_root_address_calculated
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_final_index_sum_regn_Update/$exit
      -- 
    ack_1323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_537_index_offset_ack_1, ack => convTranspose_CP_39_elements(197)); -- 
    req_1332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(197), ack => addr_of_538_final_reg_req_0); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/addr_of_538_request/ack
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/addr_of_538_request/$exit
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/addr_of_538_sample_completed_
      -- 
    ack_1333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_538_final_reg_ack_0, ack => convTranspose_CP_39_elements(198)); -- 
    -- CP-element group 199:  fork  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	521 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	255 
    -- CP-element group 199:  members (19) 
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/addr_of_538_complete/$exit
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/addr_of_538_complete/ack
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/addr_of_538_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_base_address_calculated
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_word_address_calculated
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_root_address_calculated
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_base_address_resized
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_base_addr_resize/$entry
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_base_addr_resize/$exit
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_base_addr_resize/base_resize_req
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_base_addr_resize/base_resize_ack
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_base_plus_offset/$entry
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_base_plus_offset/$exit
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_base_plus_offset/sum_rename_req
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_base_plus_offset/sum_rename_ack
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_word_addrgen/$entry
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_word_addrgen/$exit
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_word_addrgen/root_register_req
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_word_addrgen/root_register_ack
      -- 
    ack_1338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_538_final_reg_ack_1, ack => convTranspose_CP_39_elements(199)); -- 
    -- CP-element group 200:  transition  input  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	521 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (6) 
      -- CP-element group 200: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_541_update_start_
      -- CP-element group 200: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_541_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_541_Update/cr
      -- CP-element group 200: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_541_Update/$entry
      -- CP-element group 200: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_541_Sample/ra
      -- CP-element group 200: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_541_Sample/$exit
      -- 
    ra_1347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_541_inst_ack_0, ack => convTranspose_CP_39_elements(200)); -- 
    cr_1351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(200), ack => RPIPE_ConvTranspose_input_pipe_541_inst_req_1); -- 
    -- CP-element group 201:  fork  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201: 	204 
    -- CP-element group 201: 	206 
    -- CP-element group 201:  members (12) 
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_548_Sample/$entry
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_548_Sample/rr
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_548_sample_start_
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_543_Sample/$entry
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_543_sample_start_
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_541_Update/ca
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_541_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_541_update_completed_
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_543_Sample/req
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_557_sample_start_
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_557_Sample/$entry
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_557_Sample/rr
      -- 
    ca_1352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_541_inst_ack_1, ack => convTranspose_CP_39_elements(201)); -- 
    req_1360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(201), ack => WPIPE_ConvTranspose_output_pipe_543_inst_req_0); -- 
    rr_1374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(201), ack => type_cast_548_inst_req_0); -- 
    rr_1388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(201), ack => RPIPE_ConvTranspose_input_pipe_557_inst_req_0); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_543_Update/req
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_543_Sample/$exit
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_543_Sample/ack
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_543_Update/$entry
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_543_update_start_
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_543_sample_completed_
      -- 
    ack_1361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_543_inst_ack_0, ack => convTranspose_CP_39_elements(202)); -- 
    req_1365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(202), ack => WPIPE_ConvTranspose_output_pipe_543_inst_req_1); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	208 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_543_Update/$exit
      -- CP-element group 203: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_543_Update/ack
      -- CP-element group 203: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_543_update_completed_
      -- 
    ack_1366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_543_inst_ack_1, ack => convTranspose_CP_39_elements(203)); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	201 
    -- CP-element group 204: successors 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_548_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_548_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_548_Sample/ra
      -- 
    ra_1375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_548_inst_ack_0, ack => convTranspose_CP_39_elements(204)); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	521 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	255 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_548_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_548_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_548_Update/ca
      -- 
    ca_1380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_548_inst_ack_1, ack => convTranspose_CP_39_elements(205)); -- 
    -- CP-element group 206:  transition  input  output  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	201 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (6) 
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_557_sample_completed_
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_557_update_start_
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_557_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_557_Sample/ra
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_557_Update/$entry
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_557_Update/cr
      -- 
    ra_1389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_557_inst_ack_0, ack => convTranspose_CP_39_elements(206)); -- 
    cr_1393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(206), ack => RPIPE_ConvTranspose_input_pipe_557_inst_req_1); -- 
    -- CP-element group 207:  fork  transition  input  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207: 	211 
    -- CP-element group 207: 	213 
    -- CP-element group 207:  members (9) 
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_557_update_completed_
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_557_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_557_Update/ca
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_564_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_564_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_564_Sample/rr
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_578_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_578_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_578_Sample/rr
      -- 
    ca_1394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_557_inst_ack_1, ack => convTranspose_CP_39_elements(207)); -- 
    rr_1416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(207), ack => type_cast_564_inst_req_0); -- 
    rr_1430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(207), ack => RPIPE_ConvTranspose_input_pipe_578_inst_req_0); -- 
    -- CP-element group 208:  join  transition  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	203 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_559_sample_start_
      -- CP-element group 208: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_559_Sample/$entry
      -- CP-element group 208: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_559_Sample/req
      -- 
    req_1402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(208), ack => WPIPE_ConvTranspose_output_pipe_559_inst_req_0); -- 
    convTranspose_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(203) & convTranspose_CP_39_elements(207);
      gj_convTranspose_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  transition  input  output  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209:  members (6) 
      -- CP-element group 209: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_559_sample_completed_
      -- CP-element group 209: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_559_update_start_
      -- CP-element group 209: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_559_Sample/$exit
      -- CP-element group 209: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_559_Sample/ack
      -- CP-element group 209: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_559_Update/$entry
      -- CP-element group 209: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_559_Update/req
      -- 
    ack_1403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_559_inst_ack_0, ack => convTranspose_CP_39_elements(209)); -- 
    req_1407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(209), ack => WPIPE_ConvTranspose_output_pipe_559_inst_req_1); -- 
    -- CP-element group 210:  transition  input  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	215 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_559_update_completed_
      -- CP-element group 210: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_559_Update/$exit
      -- CP-element group 210: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_559_Update/ack
      -- 
    ack_1408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_559_inst_ack_1, ack => convTranspose_CP_39_elements(210)); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	207 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_564_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_564_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_564_Sample/ra
      -- 
    ra_1417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_564_inst_ack_0, ack => convTranspose_CP_39_elements(211)); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	521 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	255 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_564_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_564_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_564_Update/ca
      -- 
    ca_1422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_564_inst_ack_1, ack => convTranspose_CP_39_elements(212)); -- 
    -- CP-element group 213:  transition  input  output  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	207 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213:  members (6) 
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_578_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_578_update_start_
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_578_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_578_Sample/ra
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_578_Update/$entry
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_578_Update/cr
      -- 
    ra_1431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_578_inst_ack_0, ack => convTranspose_CP_39_elements(213)); -- 
    cr_1435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(213), ack => RPIPE_ConvTranspose_input_pipe_578_inst_req_1); -- 
    -- CP-element group 214:  fork  transition  input  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	213 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	218 
    -- CP-element group 214: 	220 
    -- CP-element group 214: 	215 
    -- CP-element group 214:  members (9) 
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_578_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_578_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_578_Update/ca
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_585_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_585_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_585_Sample/rr
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_599_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_599_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_599_Sample/rr
      -- 
    ca_1436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_578_inst_ack_1, ack => convTranspose_CP_39_elements(214)); -- 
    rr_1472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(214), ack => RPIPE_ConvTranspose_input_pipe_599_inst_req_0); -- 
    rr_1458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(214), ack => type_cast_585_inst_req_0); -- 
    -- CP-element group 215:  join  transition  output  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	210 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_580_sample_start_
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_580_Sample/$entry
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_580_Sample/req
      -- 
    req_1444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(215), ack => WPIPE_ConvTranspose_output_pipe_580_inst_req_0); -- 
    convTranspose_cp_element_group_215: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_215"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(210) & convTranspose_CP_39_elements(214);
      gj_convTranspose_cp_element_group_215 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(215), clk => clk, reset => reset); --
    end block;
    -- CP-element group 216:  transition  input  output  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (6) 
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_580_sample_completed_
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_580_update_start_
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_580_Sample/$exit
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_580_Sample/ack
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_580_Update/$entry
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_580_Update/req
      -- 
    ack_1445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_580_inst_ack_0, ack => convTranspose_CP_39_elements(216)); -- 
    req_1449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(216), ack => WPIPE_ConvTranspose_output_pipe_580_inst_req_1); -- 
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	222 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_580_update_completed_
      -- CP-element group 217: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_580_Update/$exit
      -- CP-element group 217: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_580_Update/ack
      -- 
    ack_1450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_580_inst_ack_1, ack => convTranspose_CP_39_elements(217)); -- 
    -- CP-element group 218:  transition  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	214 
    -- CP-element group 218: successors 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_585_sample_completed_
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_585_Sample/$exit
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_585_Sample/ra
      -- 
    ra_1459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_585_inst_ack_0, ack => convTranspose_CP_39_elements(218)); -- 
    -- CP-element group 219:  transition  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	521 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	255 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_585_update_completed_
      -- CP-element group 219: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_585_Update/$exit
      -- CP-element group 219: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_585_Update/ca
      -- 
    ca_1464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_585_inst_ack_1, ack => convTranspose_CP_39_elements(219)); -- 
    -- CP-element group 220:  transition  input  output  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	214 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	221 
    -- CP-element group 220:  members (6) 
      -- CP-element group 220: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_599_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_599_update_start_
      -- CP-element group 220: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_599_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_599_Sample/ra
      -- CP-element group 220: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_599_Update/$entry
      -- CP-element group 220: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_599_Update/cr
      -- 
    ra_1473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_599_inst_ack_0, ack => convTranspose_CP_39_elements(220)); -- 
    cr_1477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(220), ack => RPIPE_ConvTranspose_input_pipe_599_inst_req_1); -- 
    -- CP-element group 221:  fork  transition  input  output  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	220 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	222 
    -- CP-element group 221: 	225 
    -- CP-element group 221: 	227 
    -- CP-element group 221:  members (9) 
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_599_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_599_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_599_Update/ca
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_606_sample_start_
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_606_Sample/$entry
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_606_Sample/rr
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_620_sample_start_
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_620_Sample/$entry
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_620_Sample/rr
      -- 
    ca_1478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_599_inst_ack_1, ack => convTranspose_CP_39_elements(221)); -- 
    rr_1500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(221), ack => type_cast_606_inst_req_0); -- 
    rr_1514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(221), ack => RPIPE_ConvTranspose_input_pipe_620_inst_req_0); -- 
    -- CP-element group 222:  join  transition  output  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	221 
    -- CP-element group 222: 	217 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_601_sample_start_
      -- CP-element group 222: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_601_Sample/$entry
      -- CP-element group 222: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_601_Sample/req
      -- 
    req_1486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(222), ack => WPIPE_ConvTranspose_output_pipe_601_inst_req_0); -- 
    convTranspose_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(221) & convTranspose_CP_39_elements(217);
      gj_convTranspose_cp_element_group_222 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (6) 
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_601_sample_completed_
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_601_update_start_
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_601_Sample/$exit
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_601_Sample/ack
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_601_Update/$entry
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_601_Update/req
      -- 
    ack_1487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_601_inst_ack_0, ack => convTranspose_CP_39_elements(223)); -- 
    req_1491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(223), ack => WPIPE_ConvTranspose_output_pipe_601_inst_req_1); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	229 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_601_update_completed_
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_601_Update/$exit
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_601_Update/ack
      -- 
    ack_1492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_601_inst_ack_1, ack => convTranspose_CP_39_elements(224)); -- 
    -- CP-element group 225:  transition  input  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	221 
    -- CP-element group 225: successors 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_606_sample_completed_
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_606_Sample/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_606_Sample/ra
      -- 
    ra_1501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_606_inst_ack_0, ack => convTranspose_CP_39_elements(225)); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	521 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	255 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_606_update_completed_
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_606_Update/$exit
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_606_Update/ca
      -- 
    ca_1506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_606_inst_ack_1, ack => convTranspose_CP_39_elements(226)); -- 
    -- CP-element group 227:  transition  input  output  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	221 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (6) 
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_620_sample_completed_
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_620_update_start_
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_620_Sample/$exit
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_620_Sample/ra
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_620_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_620_Update/cr
      -- 
    ra_1515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_620_inst_ack_0, ack => convTranspose_CP_39_elements(227)); -- 
    cr_1519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(227), ack => RPIPE_ConvTranspose_input_pipe_620_inst_req_1); -- 
    -- CP-element group 228:  fork  transition  input  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	234 
    -- CP-element group 228: 	229 
    -- CP-element group 228: 	232 
    -- CP-element group 228:  members (9) 
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_620_update_completed_
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_620_Update/$exit
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_620_Update/ca
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_627_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_627_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_627_Sample/rr
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_641_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_641_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_641_Sample/rr
      -- 
    ca_1520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_620_inst_ack_1, ack => convTranspose_CP_39_elements(228)); -- 
    rr_1556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(228), ack => RPIPE_ConvTranspose_input_pipe_641_inst_req_0); -- 
    rr_1542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(228), ack => type_cast_627_inst_req_0); -- 
    -- CP-element group 229:  join  transition  output  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	224 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_622_sample_start_
      -- CP-element group 229: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_622_Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_622_Sample/req
      -- 
    req_1528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(229), ack => WPIPE_ConvTranspose_output_pipe_622_inst_req_0); -- 
    convTranspose_cp_element_group_229: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_229"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(224) & convTranspose_CP_39_elements(228);
      gj_convTranspose_cp_element_group_229 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(229), clk => clk, reset => reset); --
    end block;
    -- CP-element group 230:  transition  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	231 
    -- CP-element group 230:  members (6) 
      -- CP-element group 230: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_622_sample_completed_
      -- CP-element group 230: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_622_update_start_
      -- CP-element group 230: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_622_Sample/$exit
      -- CP-element group 230: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_622_Sample/ack
      -- CP-element group 230: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_622_Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_622_Update/req
      -- 
    ack_1529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_622_inst_ack_0, ack => convTranspose_CP_39_elements(230)); -- 
    req_1533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(230), ack => WPIPE_ConvTranspose_output_pipe_622_inst_req_1); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	236 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_622_update_completed_
      -- CP-element group 231: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_622_Update/$exit
      -- CP-element group 231: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_622_Update/ack
      -- 
    ack_1534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_622_inst_ack_1, ack => convTranspose_CP_39_elements(231)); -- 
    -- CP-element group 232:  transition  input  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	228 
    -- CP-element group 232: successors 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_627_sample_completed_
      -- CP-element group 232: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_627_Sample/$exit
      -- CP-element group 232: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_627_Sample/ra
      -- 
    ra_1543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_627_inst_ack_0, ack => convTranspose_CP_39_elements(232)); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	521 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	255 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_627_update_completed_
      -- CP-element group 233: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_627_Update/$exit
      -- CP-element group 233: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_627_Update/ca
      -- 
    ca_1548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_627_inst_ack_1, ack => convTranspose_CP_39_elements(233)); -- 
    -- CP-element group 234:  transition  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	228 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234:  members (6) 
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_641_sample_completed_
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_641_update_start_
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_641_Sample/$exit
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_641_Sample/ra
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_641_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_641_Update/cr
      -- 
    ra_1557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_641_inst_ack_0, ack => convTranspose_CP_39_elements(234)); -- 
    cr_1561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => RPIPE_ConvTranspose_input_pipe_641_inst_req_1); -- 
    -- CP-element group 235:  fork  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235: 	239 
    -- CP-element group 235: 	241 
    -- CP-element group 235:  members (9) 
      -- CP-element group 235: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_641_update_completed_
      -- CP-element group 235: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_641_Update/$exit
      -- CP-element group 235: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_641_Update/ca
      -- CP-element group 235: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_648_sample_start_
      -- CP-element group 235: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_648_Sample/$entry
      -- CP-element group 235: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_648_Sample/rr
      -- CP-element group 235: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_662_sample_start_
      -- CP-element group 235: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_662_Sample/$entry
      -- CP-element group 235: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_662_Sample/rr
      -- 
    ca_1562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_641_inst_ack_1, ack => convTranspose_CP_39_elements(235)); -- 
    rr_1584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(235), ack => type_cast_648_inst_req_0); -- 
    rr_1598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(235), ack => RPIPE_ConvTranspose_input_pipe_662_inst_req_0); -- 
    -- CP-element group 236:  join  transition  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: 	231 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_643_sample_start_
      -- CP-element group 236: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_643_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_643_Sample/req
      -- 
    req_1570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(236), ack => WPIPE_ConvTranspose_output_pipe_643_inst_req_0); -- 
    convTranspose_cp_element_group_236: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_236"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(235) & convTranspose_CP_39_elements(231);
      gj_convTranspose_cp_element_group_236 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(236), clk => clk, reset => reset); --
    end block;
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_643_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_643_update_start_
      -- CP-element group 237: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_643_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_643_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_643_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_643_Update/req
      -- 
    ack_1571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_643_inst_ack_0, ack => convTranspose_CP_39_elements(237)); -- 
    req_1575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(237), ack => WPIPE_ConvTranspose_output_pipe_643_inst_req_1); -- 
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	243 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_643_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_643_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_643_Update/ack
      -- 
    ack_1576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_643_inst_ack_1, ack => convTranspose_CP_39_elements(238)); -- 
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	235 
    -- CP-element group 239: successors 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_648_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_648_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_648_Sample/ra
      -- 
    ra_1585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_648_inst_ack_0, ack => convTranspose_CP_39_elements(239)); -- 
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	521 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	255 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_648_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_648_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_648_Update/ca
      -- 
    ca_1590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_648_inst_ack_1, ack => convTranspose_CP_39_elements(240)); -- 
    -- CP-element group 241:  transition  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	235 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_662_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_662_update_start_
      -- CP-element group 241: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_662_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_662_Sample/ra
      -- CP-element group 241: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_662_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_662_Update/cr
      -- 
    ra_1599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_662_inst_ack_0, ack => convTranspose_CP_39_elements(241)); -- 
    cr_1603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(241), ack => RPIPE_ConvTranspose_input_pipe_662_inst_req_1); -- 
    -- CP-element group 242:  fork  transition  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242: 	246 
    -- CP-element group 242: 	248 
    -- CP-element group 242:  members (9) 
      -- CP-element group 242: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_662_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_662_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_662_Update/ca
      -- CP-element group 242: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_669_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_669_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_669_Sample/rr
      -- CP-element group 242: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_683_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_683_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_683_Sample/rr
      -- 
    ca_1604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_662_inst_ack_1, ack => convTranspose_CP_39_elements(242)); -- 
    rr_1626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(242), ack => type_cast_669_inst_req_0); -- 
    rr_1640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(242), ack => RPIPE_ConvTranspose_input_pipe_683_inst_req_0); -- 
    -- CP-element group 243:  join  transition  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	238 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_664_sample_start_
      -- CP-element group 243: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_664_Sample/$entry
      -- CP-element group 243: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_664_Sample/req
      -- 
    req_1612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(243), ack => WPIPE_ConvTranspose_output_pipe_664_inst_req_0); -- 
    convTranspose_cp_element_group_243: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_243"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(238) & convTranspose_CP_39_elements(242);
      gj_convTranspose_cp_element_group_243 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(243), clk => clk, reset => reset); --
    end block;
    -- CP-element group 244:  transition  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_664_sample_completed_
      -- CP-element group 244: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_664_update_start_
      -- CP-element group 244: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_664_Sample/$exit
      -- CP-element group 244: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_664_Sample/ack
      -- CP-element group 244: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_664_Update/$entry
      -- CP-element group 244: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_664_Update/req
      -- 
    ack_1613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_664_inst_ack_0, ack => convTranspose_CP_39_elements(244)); -- 
    req_1617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(244), ack => WPIPE_ConvTranspose_output_pipe_664_inst_req_1); -- 
    -- CP-element group 245:  transition  input  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	250 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_664_update_completed_
      -- CP-element group 245: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_664_Update/$exit
      -- CP-element group 245: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_664_Update/ack
      -- 
    ack_1618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_664_inst_ack_1, ack => convTranspose_CP_39_elements(245)); -- 
    -- CP-element group 246:  transition  input  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	242 
    -- CP-element group 246: successors 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_669_sample_completed_
      -- CP-element group 246: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_669_Sample/$exit
      -- CP-element group 246: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_669_Sample/ra
      -- 
    ra_1627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_669_inst_ack_0, ack => convTranspose_CP_39_elements(246)); -- 
    -- CP-element group 247:  transition  input  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	521 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	255 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_669_update_completed_
      -- CP-element group 247: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_669_Update/$exit
      -- CP-element group 247: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_669_Update/ca
      -- 
    ca_1632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_669_inst_ack_1, ack => convTranspose_CP_39_elements(247)); -- 
    -- CP-element group 248:  transition  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	242 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (6) 
      -- CP-element group 248: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_683_sample_completed_
      -- CP-element group 248: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_683_update_start_
      -- CP-element group 248: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_683_Sample/$exit
      -- CP-element group 248: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_683_Sample/ra
      -- CP-element group 248: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_683_Update/$entry
      -- CP-element group 248: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_683_Update/cr
      -- 
    ra_1641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_683_inst_ack_0, ack => convTranspose_CP_39_elements(248)); -- 
    cr_1645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(248), ack => RPIPE_ConvTranspose_input_pipe_683_inst_req_1); -- 
    -- CP-element group 249:  fork  transition  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249: 	253 
    -- CP-element group 249:  members (6) 
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_683_update_completed_
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_683_Update/$exit
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_683_Update/ca
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_690_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_690_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_690_Sample/rr
      -- 
    ca_1646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_683_inst_ack_1, ack => convTranspose_CP_39_elements(249)); -- 
    rr_1668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(249), ack => type_cast_690_inst_req_0); -- 
    -- CP-element group 250:  join  transition  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	245 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_685_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_685_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_685_Sample/req
      -- 
    req_1654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(250), ack => WPIPE_ConvTranspose_output_pipe_685_inst_req_0); -- 
    convTranspose_cp_element_group_250: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_250"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(245) & convTranspose_CP_39_elements(249);
      gj_convTranspose_cp_element_group_250 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(250), clk => clk, reset => reset); --
    end block;
    -- CP-element group 251:  transition  input  output  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (6) 
      -- CP-element group 251: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_685_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_685_update_start_
      -- CP-element group 251: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_685_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_685_Sample/ack
      -- CP-element group 251: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_685_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_685_Update/req
      -- 
    ack_1655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_685_inst_ack_0, ack => convTranspose_CP_39_elements(251)); -- 
    req_1659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(251), ack => WPIPE_ConvTranspose_output_pipe_685_inst_req_1); -- 
    -- CP-element group 252:  transition  input  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	258 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_685_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_685_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/WPIPE_ConvTranspose_output_pipe_685_Update/ack
      -- 
    ack_1660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_685_inst_ack_1, ack => convTranspose_CP_39_elements(252)); -- 
    -- CP-element group 253:  transition  input  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	249 
    -- CP-element group 253: successors 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_690_sample_completed_
      -- CP-element group 253: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_690_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_690_Sample/ra
      -- 
    ra_1669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_690_inst_ack_0, ack => convTranspose_CP_39_elements(253)); -- 
    -- CP-element group 254:  transition  input  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	521 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_690_update_completed_
      -- CP-element group 254: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_690_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_690_Update/ca
      -- 
    ca_1674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_690_inst_ack_1, ack => convTranspose_CP_39_elements(254)); -- 
    -- CP-element group 255:  join  transition  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	199 
    -- CP-element group 255: 	205 
    -- CP-element group 255: 	240 
    -- CP-element group 255: 	247 
    -- CP-element group 255: 	219 
    -- CP-element group 255: 	254 
    -- CP-element group 255: 	226 
    -- CP-element group 255: 	233 
    -- CP-element group 255: 	212 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (9) 
      -- CP-element group 255: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_sample_start_
      -- CP-element group 255: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_Sample/$entry
      -- CP-element group 255: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_Sample/ptr_deref_698_Split/$entry
      -- CP-element group 255: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_Sample/ptr_deref_698_Split/$exit
      -- CP-element group 255: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_Sample/ptr_deref_698_Split/split_req
      -- CP-element group 255: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_Sample/ptr_deref_698_Split/split_ack
      -- CP-element group 255: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_Sample/word_access_start/$entry
      -- CP-element group 255: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_Sample/word_access_start/word_0/$entry
      -- CP-element group 255: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_Sample/word_access_start/word_0/rr
      -- 
    rr_1712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(255), ack => ptr_deref_698_store_0_req_0); -- 
    convTranspose_cp_element_group_255: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_255"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(199) & convTranspose_CP_39_elements(205) & convTranspose_CP_39_elements(240) & convTranspose_CP_39_elements(247) & convTranspose_CP_39_elements(219) & convTranspose_CP_39_elements(254) & convTranspose_CP_39_elements(226) & convTranspose_CP_39_elements(233) & convTranspose_CP_39_elements(212);
      gj_convTranspose_cp_element_group_255 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(255), clk => clk, reset => reset); --
    end block;
    -- CP-element group 256:  transition  input  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256:  members (5) 
      -- CP-element group 256: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_sample_completed_
      -- CP-element group 256: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_Sample/$exit
      -- CP-element group 256: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_Sample/word_access_start/$exit
      -- CP-element group 256: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_Sample/word_access_start/word_0/$exit
      -- CP-element group 256: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_Sample/word_access_start/word_0/ra
      -- 
    ra_1713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_698_store_0_ack_0, ack => convTranspose_CP_39_elements(256)); -- 
    -- CP-element group 257:  transition  input  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	521 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (5) 
      -- CP-element group 257: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_update_completed_
      -- CP-element group 257: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_Update/$exit
      -- CP-element group 257: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_Update/word_access_complete/$exit
      -- CP-element group 257: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_Update/word_access_complete/word_0/$exit
      -- CP-element group 257: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_Update/word_access_complete/word_0/ca
      -- 
    ca_1724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_698_store_0_ack_1, ack => convTranspose_CP_39_elements(257)); -- 
    -- CP-element group 258:  branch  join  transition  place  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	196 
    -- CP-element group 258: 	252 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258: 	260 
    -- CP-element group 258:  members (10) 
      -- CP-element group 258: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711__exit__
      -- CP-element group 258: 	 branch_block_stmt_33/if_stmt_712__entry__
      -- CP-element group 258: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/$exit
      -- CP-element group 258: 	 branch_block_stmt_33/if_stmt_712_dead_link/$entry
      -- CP-element group 258: 	 branch_block_stmt_33/if_stmt_712_eval_test/$entry
      -- CP-element group 258: 	 branch_block_stmt_33/if_stmt_712_eval_test/$exit
      -- CP-element group 258: 	 branch_block_stmt_33/if_stmt_712_eval_test/branch_req
      -- CP-element group 258: 	 branch_block_stmt_33/R_exitcond3_713_place
      -- CP-element group 258: 	 branch_block_stmt_33/if_stmt_712_if_link/$entry
      -- CP-element group 258: 	 branch_block_stmt_33/if_stmt_712_else_link/$entry
      -- 
    branch_req_1732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(258), ack => if_stmt_712_branch_req_0); -- 
    convTranspose_cp_element_group_258: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_258"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(196) & convTranspose_CP_39_elements(252) & convTranspose_CP_39_elements(257);
      gj_convTranspose_cp_element_group_258 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(258), clk => clk, reset => reset); --
    end block;
    -- CP-element group 259:  merge  transition  place  input  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	515 
    -- CP-element group 259:  members (13) 
      -- CP-element group 259: 	 branch_block_stmt_33/merge_stmt_472__exit__
      -- CP-element group 259: 	 branch_block_stmt_33/forx_xcond302x_xpreheaderx_xloopexit_forx_xcond302x_xpreheader
      -- CP-element group 259: 	 branch_block_stmt_33/if_stmt_712_if_link/$exit
      -- CP-element group 259: 	 branch_block_stmt_33/if_stmt_712_if_link/if_choice_transition
      -- CP-element group 259: 	 branch_block_stmt_33/forx_xbody_forx_xcond302x_xpreheaderx_xloopexit
      -- CP-element group 259: 	 branch_block_stmt_33/forx_xbody_forx_xcond302x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 259: 	 branch_block_stmt_33/forx_xbody_forx_xcond302x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 259: 	 branch_block_stmt_33/merge_stmt_472_PhiReqMerge
      -- CP-element group 259: 	 branch_block_stmt_33/merge_stmt_472_PhiAck/$entry
      -- CP-element group 259: 	 branch_block_stmt_33/merge_stmt_472_PhiAck/$exit
      -- CP-element group 259: 	 branch_block_stmt_33/merge_stmt_472_PhiAck/dummy
      -- CP-element group 259: 	 branch_block_stmt_33/forx_xcond302x_xpreheaderx_xloopexit_forx_xcond302x_xpreheader_PhiReq/$entry
      -- CP-element group 259: 	 branch_block_stmt_33/forx_xcond302x_xpreheaderx_xloopexit_forx_xcond302x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_712_branch_ack_1, ack => convTranspose_CP_39_elements(259)); -- 
    -- CP-element group 260:  fork  transition  place  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	517 
    -- CP-element group 260: 	518 
    -- CP-element group 260:  members (12) 
      -- CP-element group 260: 	 branch_block_stmt_33/if_stmt_712_else_link/$exit
      -- CP-element group 260: 	 branch_block_stmt_33/if_stmt_712_else_link/else_choice_transition
      -- CP-element group 260: 	 branch_block_stmt_33/forx_xbody_forx_xbody
      -- CP-element group 260: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 260: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_525/$entry
      -- CP-element group 260: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_525/phi_stmt_525_sources/$entry
      -- CP-element group 260: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_525/phi_stmt_525_sources/type_cast_531/$entry
      -- CP-element group 260: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_525/phi_stmt_525_sources/type_cast_531/SplitProtocol/$entry
      -- CP-element group 260: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_525/phi_stmt_525_sources/type_cast_531/SplitProtocol/Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_525/phi_stmt_525_sources/type_cast_531/SplitProtocol/Sample/rr
      -- CP-element group 260: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_525/phi_stmt_525_sources/type_cast_531/SplitProtocol/Update/$entry
      -- CP-element group 260: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_525/phi_stmt_525_sources/type_cast_531/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_712_branch_ack_0, ack => convTranspose_CP_39_elements(260)); -- 
    rr_3660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(260), ack => type_cast_531_inst_req_0); -- 
    cr_3665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(260), ack => type_cast_531_inst_req_1); -- 
    -- CP-element group 261:  transition  input  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	192 
    -- CP-element group 261: successors 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_724_to_assign_stmt_753/type_cast_739_sample_completed_
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_724_to_assign_stmt_753/type_cast_739_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_724_to_assign_stmt_753/type_cast_739_Sample/ra
      -- 
    ra_1755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_739_inst_ack_0, ack => convTranspose_CP_39_elements(261)); -- 
    -- CP-element group 262:  transition  place  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	192 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	522 
    -- CP-element group 262:  members (9) 
      -- CP-element group 262: 	 branch_block_stmt_33/assign_stmt_724_to_assign_stmt_753__exit__
      -- CP-element group 262: 	 branch_block_stmt_33/bbx_xnph573_forx_xbody308
      -- CP-element group 262: 	 branch_block_stmt_33/assign_stmt_724_to_assign_stmt_753/$exit
      -- CP-element group 262: 	 branch_block_stmt_33/assign_stmt_724_to_assign_stmt_753/type_cast_739_update_completed_
      -- CP-element group 262: 	 branch_block_stmt_33/assign_stmt_724_to_assign_stmt_753/type_cast_739_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_33/assign_stmt_724_to_assign_stmt_753/type_cast_739_Update/ca
      -- CP-element group 262: 	 branch_block_stmt_33/bbx_xnph573_forx_xbody308_PhiReq/$entry
      -- CP-element group 262: 	 branch_block_stmt_33/bbx_xnph573_forx_xbody308_PhiReq/phi_stmt_756/$entry
      -- CP-element group 262: 	 branch_block_stmt_33/bbx_xnph573_forx_xbody308_PhiReq/phi_stmt_756/phi_stmt_756_sources/$entry
      -- 
    ca_1760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_739_inst_ack_1, ack => convTranspose_CP_39_elements(262)); -- 
    -- CP-element group 263:  transition  input  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	527 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	325 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_final_index_sum_regn_sample_complete
      -- CP-element group 263: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_final_index_sum_regn_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_final_index_sum_regn_Sample/ack
      -- 
    ack_1789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_768_index_offset_ack_0, ack => convTranspose_CP_39_elements(263)); -- 
    -- CP-element group 264:  transition  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	527 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (11) 
      -- CP-element group 264: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/addr_of_769_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_root_address_calculated
      -- CP-element group 264: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_offset_calculated
      -- CP-element group 264: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_final_index_sum_regn_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_final_index_sum_regn_Update/ack
      -- CP-element group 264: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_base_plus_offset/$entry
      -- CP-element group 264: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_base_plus_offset/$exit
      -- CP-element group 264: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_base_plus_offset/sum_rename_req
      -- CP-element group 264: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_base_plus_offset/sum_rename_ack
      -- CP-element group 264: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/addr_of_769_request/$entry
      -- CP-element group 264: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/addr_of_769_request/req
      -- 
    ack_1794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_768_index_offset_ack_1, ack => convTranspose_CP_39_elements(264)); -- 
    req_1803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(264), ack => addr_of_769_final_reg_req_0); -- 
    -- CP-element group 265:  transition  input  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/addr_of_769_sample_completed_
      -- CP-element group 265: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/addr_of_769_request/$exit
      -- CP-element group 265: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/addr_of_769_request/ack
      -- 
    ack_1804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_769_final_reg_ack_0, ack => convTranspose_CP_39_elements(265)); -- 
    -- CP-element group 266:  fork  transition  input  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	527 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	322 
    -- CP-element group 266:  members (19) 
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_word_addrgen/root_register_ack
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_word_addrgen/root_register_req
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_word_addrgen/$exit
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_word_addrgen/$entry
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_base_plus_offset/sum_rename_ack
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_base_plus_offset/sum_rename_req
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_base_plus_offset/$exit
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_base_plus_offset/$entry
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_base_addr_resize/base_resize_ack
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_base_addr_resize/base_resize_req
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_base_addr_resize/$exit
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_base_addr_resize/$entry
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_base_address_resized
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_root_address_calculated
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_word_address_calculated
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_base_address_calculated
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/addr_of_769_update_completed_
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/addr_of_769_complete/$exit
      -- CP-element group 266: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/addr_of_769_complete/ack
      -- 
    ack_1809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_769_final_reg_ack_1, ack => convTranspose_CP_39_elements(266)); -- 
    -- CP-element group 267:  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	527 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (6) 
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_772_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_772_update_start_
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_772_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_772_Sample/ra
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_772_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_772_Update/cr
      -- 
    ra_1818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_772_inst_ack_0, ack => convTranspose_CP_39_elements(267)); -- 
    cr_1822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(267), ack => RPIPE_ConvTranspose_input_pipe_772_inst_req_1); -- 
    -- CP-element group 268:  fork  transition  input  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268: 	271 
    -- CP-element group 268: 	273 
    -- CP-element group 268:  members (12) 
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_772_update_completed_
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_772_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_772_Update/ca
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_774_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_774_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_774_Sample/req
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_779_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_779_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_779_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_788_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_788_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_788_Sample/rr
      -- 
    ca_1823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_772_inst_ack_1, ack => convTranspose_CP_39_elements(268)); -- 
    req_1831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(268), ack => WPIPE_ConvTranspose_output_pipe_774_inst_req_0); -- 
    rr_1845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(268), ack => type_cast_779_inst_req_0); -- 
    rr_1859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(268), ack => RPIPE_ConvTranspose_input_pipe_788_inst_req_0); -- 
    -- CP-element group 269:  transition  input  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (6) 
      -- CP-element group 269: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_774_sample_completed_
      -- CP-element group 269: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_774_update_start_
      -- CP-element group 269: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_774_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_774_Sample/ack
      -- CP-element group 269: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_774_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_774_Update/req
      -- 
    ack_1832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_774_inst_ack_0, ack => convTranspose_CP_39_elements(269)); -- 
    req_1836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(269), ack => WPIPE_ConvTranspose_output_pipe_774_inst_req_1); -- 
    -- CP-element group 270:  transition  input  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	275 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_774_update_completed_
      -- CP-element group 270: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_774_Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_774_Update/ack
      -- 
    ack_1837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_774_inst_ack_1, ack => convTranspose_CP_39_elements(270)); -- 
    -- CP-element group 271:  transition  input  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	268 
    -- CP-element group 271: successors 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_779_sample_completed_
      -- CP-element group 271: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_779_Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_779_Sample/ra
      -- 
    ra_1846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_779_inst_ack_0, ack => convTranspose_CP_39_elements(271)); -- 
    -- CP-element group 272:  transition  input  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	527 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	322 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_779_update_completed_
      -- CP-element group 272: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_779_Update/$exit
      -- CP-element group 272: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_779_Update/ca
      -- 
    ca_1851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_779_inst_ack_1, ack => convTranspose_CP_39_elements(272)); -- 
    -- CP-element group 273:  transition  input  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	268 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (6) 
      -- CP-element group 273: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_788_sample_completed_
      -- CP-element group 273: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_788_update_start_
      -- CP-element group 273: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_788_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_788_Sample/ra
      -- CP-element group 273: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_788_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_788_Update/cr
      -- 
    ra_1860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_788_inst_ack_0, ack => convTranspose_CP_39_elements(273)); -- 
    cr_1864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(273), ack => RPIPE_ConvTranspose_input_pipe_788_inst_req_1); -- 
    -- CP-element group 274:  fork  transition  input  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274: 	278 
    -- CP-element group 274: 	280 
    -- CP-element group 274:  members (9) 
      -- CP-element group 274: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_788_update_completed_
      -- CP-element group 274: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_788_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_788_Update/ca
      -- CP-element group 274: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_795_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_795_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_795_Sample/rr
      -- CP-element group 274: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_809_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_809_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_809_Sample/rr
      -- 
    ca_1865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_788_inst_ack_1, ack => convTranspose_CP_39_elements(274)); -- 
    rr_1887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(274), ack => type_cast_795_inst_req_0); -- 
    rr_1901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(274), ack => RPIPE_ConvTranspose_input_pipe_809_inst_req_0); -- 
    -- CP-element group 275:  join  transition  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	270 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_790_sample_start_
      -- CP-element group 275: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_790_Sample/$entry
      -- CP-element group 275: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_790_Sample/req
      -- 
    req_1873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(275), ack => WPIPE_ConvTranspose_output_pipe_790_inst_req_0); -- 
    convTranspose_cp_element_group_275: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_275"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(270) & convTranspose_CP_39_elements(274);
      gj_convTranspose_cp_element_group_275 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(275), clk => clk, reset => reset); --
    end block;
    -- CP-element group 276:  transition  input  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (6) 
      -- CP-element group 276: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_790_sample_completed_
      -- CP-element group 276: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_790_update_start_
      -- CP-element group 276: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_790_Sample/$exit
      -- CP-element group 276: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_790_Sample/ack
      -- CP-element group 276: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_790_Update/$entry
      -- CP-element group 276: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_790_Update/req
      -- 
    ack_1874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_790_inst_ack_0, ack => convTranspose_CP_39_elements(276)); -- 
    req_1878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(276), ack => WPIPE_ConvTranspose_output_pipe_790_inst_req_1); -- 
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	282 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_790_update_completed_
      -- CP-element group 277: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_790_Update/$exit
      -- CP-element group 277: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_790_Update/ack
      -- 
    ack_1879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_790_inst_ack_1, ack => convTranspose_CP_39_elements(277)); -- 
    -- CP-element group 278:  transition  input  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	274 
    -- CP-element group 278: successors 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_795_sample_completed_
      -- CP-element group 278: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_795_Sample/$exit
      -- CP-element group 278: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_795_Sample/ra
      -- 
    ra_1888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_795_inst_ack_0, ack => convTranspose_CP_39_elements(278)); -- 
    -- CP-element group 279:  transition  input  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	527 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	322 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_795_update_completed_
      -- CP-element group 279: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_795_Update/$exit
      -- CP-element group 279: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_795_Update/ca
      -- 
    ca_1893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_795_inst_ack_1, ack => convTranspose_CP_39_elements(279)); -- 
    -- CP-element group 280:  transition  input  output  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	274 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280:  members (6) 
      -- CP-element group 280: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_809_sample_completed_
      -- CP-element group 280: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_809_update_start_
      -- CP-element group 280: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_809_Sample/$exit
      -- CP-element group 280: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_809_Sample/ra
      -- CP-element group 280: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_809_Update/$entry
      -- CP-element group 280: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_809_Update/cr
      -- 
    ra_1902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_809_inst_ack_0, ack => convTranspose_CP_39_elements(280)); -- 
    cr_1906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(280), ack => RPIPE_ConvTranspose_input_pipe_809_inst_req_1); -- 
    -- CP-element group 281:  fork  transition  input  output  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	282 
    -- CP-element group 281: 	285 
    -- CP-element group 281: 	287 
    -- CP-element group 281:  members (9) 
      -- CP-element group 281: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_816_Sample/$entry
      -- CP-element group 281: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_816_Sample/rr
      -- CP-element group 281: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_816_sample_start_
      -- CP-element group 281: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_830_Sample/$entry
      -- CP-element group 281: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_830_Sample/rr
      -- CP-element group 281: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_830_sample_start_
      -- CP-element group 281: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_809_update_completed_
      -- CP-element group 281: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_809_Update/$exit
      -- CP-element group 281: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_809_Update/ca
      -- 
    ca_1907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_809_inst_ack_1, ack => convTranspose_CP_39_elements(281)); -- 
    rr_1929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(281), ack => type_cast_816_inst_req_0); -- 
    rr_1943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(281), ack => RPIPE_ConvTranspose_input_pipe_830_inst_req_0); -- 
    -- CP-element group 282:  join  transition  output  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	277 
    -- CP-element group 282: 	281 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_811_sample_start_
      -- CP-element group 282: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_811_Sample/$entry
      -- CP-element group 282: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_811_Sample/req
      -- 
    req_1915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(282), ack => WPIPE_ConvTranspose_output_pipe_811_inst_req_0); -- 
    convTranspose_cp_element_group_282: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_282"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(277) & convTranspose_CP_39_elements(281);
      gj_convTranspose_cp_element_group_282 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(282), clk => clk, reset => reset); --
    end block;
    -- CP-element group 283:  transition  input  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (6) 
      -- CP-element group 283: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_811_Update/req
      -- CP-element group 283: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_811_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_811_sample_completed_
      -- CP-element group 283: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_811_update_start_
      -- CP-element group 283: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_811_Sample/$exit
      -- CP-element group 283: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_811_Sample/ack
      -- 
    ack_1916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_811_inst_ack_0, ack => convTranspose_CP_39_elements(283)); -- 
    req_1920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(283), ack => WPIPE_ConvTranspose_output_pipe_811_inst_req_1); -- 
    -- CP-element group 284:  transition  input  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	289 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_811_Update/ack
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_811_Update/$exit
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_811_update_completed_
      -- 
    ack_1921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_811_inst_ack_1, ack => convTranspose_CP_39_elements(284)); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	281 
    -- CP-element group 285: successors 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_816_sample_completed_
      -- CP-element group 285: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_816_Sample/$exit
      -- CP-element group 285: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_816_Sample/ra
      -- 
    ra_1930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_816_inst_ack_0, ack => convTranspose_CP_39_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	527 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	322 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_816_Update/$exit
      -- CP-element group 286: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_816_Update/ca
      -- CP-element group 286: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_816_update_completed_
      -- 
    ca_1935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_816_inst_ack_1, ack => convTranspose_CP_39_elements(286)); -- 
    -- CP-element group 287:  transition  input  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	281 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (6) 
      -- CP-element group 287: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_830_Sample/$exit
      -- CP-element group 287: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_830_Sample/ra
      -- CP-element group 287: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_830_Update/cr
      -- CP-element group 287: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_830_sample_completed_
      -- CP-element group 287: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_830_update_start_
      -- CP-element group 287: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_830_Update/$entry
      -- 
    ra_1944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_830_inst_ack_0, ack => convTranspose_CP_39_elements(287)); -- 
    cr_1948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(287), ack => RPIPE_ConvTranspose_input_pipe_830_inst_req_1); -- 
    -- CP-element group 288:  fork  transition  input  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288: 	292 
    -- CP-element group 288: 	294 
    -- CP-element group 288:  members (9) 
      -- CP-element group 288: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_851_Sample/rr
      -- CP-element group 288: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_830_update_completed_
      -- CP-element group 288: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_830_Update/$exit
      -- CP-element group 288: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_830_Update/ca
      -- CP-element group 288: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_851_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_851_sample_start_
      -- CP-element group 288: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_837_Sample/rr
      -- CP-element group 288: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_837_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_837_sample_start_
      -- 
    ca_1949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_830_inst_ack_1, ack => convTranspose_CP_39_elements(288)); -- 
    rr_1971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(288), ack => type_cast_837_inst_req_0); -- 
    rr_1985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(288), ack => RPIPE_ConvTranspose_input_pipe_851_inst_req_0); -- 
    -- CP-element group 289:  join  transition  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	284 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_832_sample_start_
      -- CP-element group 289: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_832_Sample/req
      -- CP-element group 289: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_832_Sample/$entry
      -- 
    req_1957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(289), ack => WPIPE_ConvTranspose_output_pipe_832_inst_req_0); -- 
    convTranspose_cp_element_group_289: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_289"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(284) & convTranspose_CP_39_elements(288);
      gj_convTranspose_cp_element_group_289 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(289), clk => clk, reset => reset); --
    end block;
    -- CP-element group 290:  transition  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (6) 
      -- CP-element group 290: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_832_sample_completed_
      -- CP-element group 290: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_832_update_start_
      -- CP-element group 290: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_832_Update/req
      -- CP-element group 290: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_832_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_832_Sample/ack
      -- CP-element group 290: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_832_Sample/$exit
      -- 
    ack_1958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_832_inst_ack_0, ack => convTranspose_CP_39_elements(290)); -- 
    req_1962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(290), ack => WPIPE_ConvTranspose_output_pipe_832_inst_req_1); -- 
    -- CP-element group 291:  transition  input  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	296 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_832_update_completed_
      -- CP-element group 291: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_832_Update/ack
      -- CP-element group 291: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_832_Update/$exit
      -- 
    ack_1963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_832_inst_ack_1, ack => convTranspose_CP_39_elements(291)); -- 
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	288 
    -- CP-element group 292: successors 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_837_Sample/ra
      -- CP-element group 292: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_837_Sample/$exit
      -- CP-element group 292: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_837_sample_completed_
      -- 
    ra_1972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_837_inst_ack_0, ack => convTranspose_CP_39_elements(292)); -- 
    -- CP-element group 293:  transition  input  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	527 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	322 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_837_Update/ca
      -- CP-element group 293: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_837_Update/$exit
      -- CP-element group 293: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_837_update_completed_
      -- 
    ca_1977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_837_inst_ack_1, ack => convTranspose_CP_39_elements(293)); -- 
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	288 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_851_Sample/$exit
      -- CP-element group 294: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_851_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_851_Update/cr
      -- CP-element group 294: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_851_Sample/ra
      -- CP-element group 294: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_851_update_start_
      -- CP-element group 294: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_851_sample_completed_
      -- 
    ra_1986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_851_inst_ack_0, ack => convTranspose_CP_39_elements(294)); -- 
    cr_1990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(294), ack => RPIPE_ConvTranspose_input_pipe_851_inst_req_1); -- 
    -- CP-element group 295:  fork  transition  input  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295: 	299 
    -- CP-element group 295: 	301 
    -- CP-element group 295:  members (9) 
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_872_Sample/rr
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_851_Update/$exit
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_858_Sample/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_858_Sample/rr
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_858_sample_start_
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_851_Update/ca
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_872_sample_start_
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_851_update_completed_
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_872_Sample/$entry
      -- 
    ca_1991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_851_inst_ack_1, ack => convTranspose_CP_39_elements(295)); -- 
    rr_2013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(295), ack => type_cast_858_inst_req_0); -- 
    rr_2027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(295), ack => RPIPE_ConvTranspose_input_pipe_872_inst_req_0); -- 
    -- CP-element group 296:  join  transition  output  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: 	291 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_853_sample_start_
      -- CP-element group 296: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_853_Sample/$entry
      -- CP-element group 296: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_853_Sample/req
      -- 
    req_1999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(296), ack => WPIPE_ConvTranspose_output_pipe_853_inst_req_0); -- 
    convTranspose_cp_element_group_296: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_296"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(295) & convTranspose_CP_39_elements(291);
      gj_convTranspose_cp_element_group_296 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(296), clk => clk, reset => reset); --
    end block;
    -- CP-element group 297:  transition  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	296 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (6) 
      -- CP-element group 297: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_853_Update/req
      -- CP-element group 297: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_853_sample_completed_
      -- CP-element group 297: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_853_Sample/ack
      -- CP-element group 297: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_853_Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_853_update_start_
      -- CP-element group 297: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_853_Sample/$exit
      -- 
    ack_2000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_853_inst_ack_0, ack => convTranspose_CP_39_elements(297)); -- 
    req_2004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(297), ack => WPIPE_ConvTranspose_output_pipe_853_inst_req_1); -- 
    -- CP-element group 298:  transition  input  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	303 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_853_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_853_update_completed_
      -- CP-element group 298: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_853_Update/ack
      -- 
    ack_2005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_853_inst_ack_1, ack => convTranspose_CP_39_elements(298)); -- 
    -- CP-element group 299:  transition  input  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	295 
    -- CP-element group 299: successors 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_858_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_858_Sample/ra
      -- CP-element group 299: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_858_sample_completed_
      -- 
    ra_2014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_858_inst_ack_0, ack => convTranspose_CP_39_elements(299)); -- 
    -- CP-element group 300:  transition  input  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	527 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	322 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_858_update_completed_
      -- CP-element group 300: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_858_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_858_Update/ca
      -- 
    ca_2019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_858_inst_ack_1, ack => convTranspose_CP_39_elements(300)); -- 
    -- CP-element group 301:  transition  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	295 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (6) 
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_872_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_872_Sample/ra
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_872_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_872_sample_completed_
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_872_Sample/$exit
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_872_update_start_
      -- 
    ra_2028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_872_inst_ack_0, ack => convTranspose_CP_39_elements(301)); -- 
    cr_2032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(301), ack => RPIPE_ConvTranspose_input_pipe_872_inst_req_1); -- 
    -- CP-element group 302:  fork  transition  input  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302: 	306 
    -- CP-element group 302: 	308 
    -- CP-element group 302:  members (9) 
      -- CP-element group 302: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_872_Update/ca
      -- CP-element group 302: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_872_Update/$exit
      -- CP-element group 302: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_893_Sample/rr
      -- CP-element group 302: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_893_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_893_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_872_update_completed_
      -- CP-element group 302: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_879_Sample/rr
      -- CP-element group 302: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_879_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_879_sample_start_
      -- 
    ca_2033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_872_inst_ack_1, ack => convTranspose_CP_39_elements(302)); -- 
    rr_2055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(302), ack => type_cast_879_inst_req_0); -- 
    rr_2069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(302), ack => RPIPE_ConvTranspose_input_pipe_893_inst_req_0); -- 
    -- CP-element group 303:  join  transition  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	298 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_874_sample_start_
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_874_Sample/req
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_874_Sample/$entry
      -- 
    req_2041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(303), ack => WPIPE_ConvTranspose_output_pipe_874_inst_req_0); -- 
    convTranspose_cp_element_group_303: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_303"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(298) & convTranspose_CP_39_elements(302);
      gj_convTranspose_cp_element_group_303 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(303), clk => clk, reset => reset); --
    end block;
    -- CP-element group 304:  transition  input  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (6) 
      -- CP-element group 304: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_874_sample_completed_
      -- CP-element group 304: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_874_update_start_
      -- CP-element group 304: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_874_Sample/$exit
      -- CP-element group 304: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_874_Sample/ack
      -- CP-element group 304: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_874_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_874_Update/req
      -- 
    ack_2042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_874_inst_ack_0, ack => convTranspose_CP_39_elements(304)); -- 
    req_2046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(304), ack => WPIPE_ConvTranspose_output_pipe_874_inst_req_1); -- 
    -- CP-element group 305:  transition  input  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	310 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_874_update_completed_
      -- CP-element group 305: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_874_Update/ack
      -- CP-element group 305: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_874_Update/$exit
      -- 
    ack_2047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_874_inst_ack_1, ack => convTranspose_CP_39_elements(305)); -- 
    -- CP-element group 306:  transition  input  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	302 
    -- CP-element group 306: successors 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_879_Sample/ra
      -- CP-element group 306: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_879_Sample/$exit
      -- CP-element group 306: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_879_sample_completed_
      -- 
    ra_2056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_879_inst_ack_0, ack => convTranspose_CP_39_elements(306)); -- 
    -- CP-element group 307:  transition  input  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	527 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	322 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_879_Update/ca
      -- CP-element group 307: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_879_Update/$exit
      -- CP-element group 307: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_879_update_completed_
      -- 
    ca_2061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_879_inst_ack_1, ack => convTranspose_CP_39_elements(307)); -- 
    -- CP-element group 308:  transition  input  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	302 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (6) 
      -- CP-element group 308: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_893_Update/cr
      -- CP-element group 308: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_893_Update/$entry
      -- CP-element group 308: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_893_Sample/ra
      -- CP-element group 308: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_893_Sample/$exit
      -- CP-element group 308: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_893_update_start_
      -- CP-element group 308: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_893_sample_completed_
      -- 
    ra_2070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_893_inst_ack_0, ack => convTranspose_CP_39_elements(308)); -- 
    cr_2074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(308), ack => RPIPE_ConvTranspose_input_pipe_893_inst_req_1); -- 
    -- CP-element group 309:  fork  transition  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309: 	313 
    -- CP-element group 309: 	315 
    -- CP-element group 309:  members (9) 
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_900_Sample/rr
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_914_Sample/$entry
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_900_Sample/$entry
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_900_sample_start_
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_914_sample_start_
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_914_Sample/rr
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_893_Update/ca
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_893_Update/$exit
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_893_update_completed_
      -- 
    ca_2075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_893_inst_ack_1, ack => convTranspose_CP_39_elements(309)); -- 
    rr_2097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(309), ack => type_cast_900_inst_req_0); -- 
    rr_2111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(309), ack => RPIPE_ConvTranspose_input_pipe_914_inst_req_0); -- 
    -- CP-element group 310:  join  transition  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	305 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_895_Sample/req
      -- CP-element group 310: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_895_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_895_sample_start_
      -- 
    req_2083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(310), ack => WPIPE_ConvTranspose_output_pipe_895_inst_req_0); -- 
    convTranspose_cp_element_group_310: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_310"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(305) & convTranspose_CP_39_elements(309);
      gj_convTranspose_cp_element_group_310 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(310), clk => clk, reset => reset); --
    end block;
    -- CP-element group 311:  transition  input  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (6) 
      -- CP-element group 311: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_895_Sample/ack
      -- CP-element group 311: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_895_Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_895_Update/req
      -- CP-element group 311: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_895_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_895_update_start_
      -- CP-element group 311: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_895_sample_completed_
      -- 
    ack_2084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_895_inst_ack_0, ack => convTranspose_CP_39_elements(311)); -- 
    req_2088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(311), ack => WPIPE_ConvTranspose_output_pipe_895_inst_req_1); -- 
    -- CP-element group 312:  transition  input  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	317 
    -- CP-element group 312:  members (3) 
      -- CP-element group 312: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_895_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_895_Update/ack
      -- CP-element group 312: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_895_update_completed_
      -- 
    ack_2089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_895_inst_ack_1, ack => convTranspose_CP_39_elements(312)); -- 
    -- CP-element group 313:  transition  input  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	309 
    -- CP-element group 313: successors 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_900_sample_completed_
      -- CP-element group 313: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_900_Sample/ra
      -- CP-element group 313: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_900_Sample/$exit
      -- 
    ra_2098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_900_inst_ack_0, ack => convTranspose_CP_39_elements(313)); -- 
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	527 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	322 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_900_update_completed_
      -- CP-element group 314: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_900_Update/$exit
      -- CP-element group 314: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_900_Update/ca
      -- 
    ca_2103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_900_inst_ack_1, ack => convTranspose_CP_39_elements(314)); -- 
    -- CP-element group 315:  transition  input  output  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	309 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	316 
    -- CP-element group 315:  members (6) 
      -- CP-element group 315: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_914_Sample/ra
      -- CP-element group 315: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_914_Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_914_Update/$entry
      -- CP-element group 315: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_914_Update/cr
      -- CP-element group 315: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_914_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_914_update_start_
      -- 
    ra_2112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_914_inst_ack_0, ack => convTranspose_CP_39_elements(315)); -- 
    cr_2116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(315), ack => RPIPE_ConvTranspose_input_pipe_914_inst_req_1); -- 
    -- CP-element group 316:  fork  transition  input  output  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	315 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316: 	320 
    -- CP-element group 316:  members (6) 
      -- CP-element group 316: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_914_Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_914_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_921_sample_start_
      -- CP-element group 316: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_914_Update/ca
      -- CP-element group 316: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_921_Sample/$entry
      -- CP-element group 316: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_921_Sample/rr
      -- 
    ca_2117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_914_inst_ack_1, ack => convTranspose_CP_39_elements(316)); -- 
    rr_2139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(316), ack => type_cast_921_inst_req_0); -- 
    -- CP-element group 317:  join  transition  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	312 
    -- CP-element group 317: 	316 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_916_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_916_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_916_Sample/req
      -- 
    req_2125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(317), ack => WPIPE_ConvTranspose_output_pipe_916_inst_req_0); -- 
    convTranspose_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(312) & convTranspose_CP_39_elements(316);
      gj_convTranspose_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  transition  input  output  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (6) 
      -- CP-element group 318: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_916_Update/$entry
      -- CP-element group 318: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_916_Update/req
      -- CP-element group 318: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_916_sample_completed_
      -- CP-element group 318: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_916_update_start_
      -- CP-element group 318: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_916_Sample/$exit
      -- CP-element group 318: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_916_Sample/ack
      -- 
    ack_2126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_916_inst_ack_0, ack => convTranspose_CP_39_elements(318)); -- 
    req_2130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(318), ack => WPIPE_ConvTranspose_output_pipe_916_inst_req_1); -- 
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	325 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_916_Update/$exit
      -- CP-element group 319: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_916_Update/ack
      -- CP-element group 319: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/WPIPE_ConvTranspose_output_pipe_916_update_completed_
      -- 
    ack_2131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_916_inst_ack_1, ack => convTranspose_CP_39_elements(319)); -- 
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	316 
    -- CP-element group 320: successors 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_921_Sample/ra
      -- CP-element group 320: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_921_sample_completed_
      -- CP-element group 320: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_921_Sample/$exit
      -- 
    ra_2140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_921_inst_ack_0, ack => convTranspose_CP_39_elements(320)); -- 
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	527 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_921_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_921_update_completed_
      -- CP-element group 321: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_921_Update/ca
      -- 
    ca_2145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_921_inst_ack_1, ack => convTranspose_CP_39_elements(321)); -- 
    -- CP-element group 322:  join  transition  output  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	300 
    -- CP-element group 322: 	307 
    -- CP-element group 322: 	314 
    -- CP-element group 322: 	321 
    -- CP-element group 322: 	266 
    -- CP-element group 322: 	272 
    -- CP-element group 322: 	279 
    -- CP-element group 322: 	286 
    -- CP-element group 322: 	293 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (9) 
      -- CP-element group 322: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_Sample/word_access_start/word_0/rr
      -- CP-element group 322: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_Sample/word_access_start/word_0/$entry
      -- CP-element group 322: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_Sample/word_access_start/$entry
      -- CP-element group 322: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_Sample/ptr_deref_929_Split/split_ack
      -- CP-element group 322: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_Sample/ptr_deref_929_Split/split_req
      -- CP-element group 322: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_Sample/ptr_deref_929_Split/$exit
      -- CP-element group 322: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_Sample/ptr_deref_929_Split/$entry
      -- CP-element group 322: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_sample_start_
      -- 
    rr_2183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(322), ack => ptr_deref_929_store_0_req_0); -- 
    convTranspose_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(300) & convTranspose_CP_39_elements(307) & convTranspose_CP_39_elements(314) & convTranspose_CP_39_elements(321) & convTranspose_CP_39_elements(266) & convTranspose_CP_39_elements(272) & convTranspose_CP_39_elements(279) & convTranspose_CP_39_elements(286) & convTranspose_CP_39_elements(293);
      gj_convTranspose_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  transition  input  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323:  members (5) 
      -- CP-element group 323: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_Sample/word_access_start/word_0/ra
      -- CP-element group 323: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_Sample/word_access_start/word_0/$exit
      -- CP-element group 323: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_Sample/word_access_start/$exit
      -- CP-element group 323: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_sample_completed_
      -- 
    ra_2184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_929_store_0_ack_0, ack => convTranspose_CP_39_elements(323)); -- 
    -- CP-element group 324:  transition  input  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	527 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (5) 
      -- CP-element group 324: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_Update/word_access_complete/word_0/$exit
      -- CP-element group 324: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_Update/word_access_complete/word_0/ca
      -- CP-element group 324: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_Update/word_access_complete/$exit
      -- CP-element group 324: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_update_completed_
      -- 
    ca_2195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_929_store_0_ack_1, ack => convTranspose_CP_39_elements(324)); -- 
    -- CP-element group 325:  branch  join  transition  place  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	319 
    -- CP-element group 325: 	324 
    -- CP-element group 325: 	263 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325: 	327 
    -- CP-element group 325:  members (10) 
      -- CP-element group 325: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942__exit__
      -- CP-element group 325: 	 branch_block_stmt_33/if_stmt_943__entry__
      -- CP-element group 325: 	 branch_block_stmt_33/if_stmt_943_eval_test/$entry
      -- CP-element group 325: 	 branch_block_stmt_33/if_stmt_943_dead_link/$entry
      -- CP-element group 325: 	 branch_block_stmt_33/if_stmt_943_eval_test/$exit
      -- CP-element group 325: 	 branch_block_stmt_33/if_stmt_943_eval_test/branch_req
      -- CP-element group 325: 	 branch_block_stmt_33/if_stmt_943_else_link/$entry
      -- CP-element group 325: 	 branch_block_stmt_33/if_stmt_943_if_link/$entry
      -- CP-element group 325: 	 branch_block_stmt_33/R_exitcond2_944_place
      -- CP-element group 325: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/$exit
      -- 
    branch_req_2203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(325), ack => if_stmt_943_branch_req_0); -- 
    convTranspose_cp_element_group_325: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_325"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(319) & convTranspose_CP_39_elements(324) & convTranspose_CP_39_elements(263);
      gj_convTranspose_cp_element_group_325 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(325), clk => clk, reset => reset); --
    end block;
    -- CP-element group 326:  merge  transition  place  input  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	528 
    -- CP-element group 326:  members (13) 
      -- CP-element group 326: 	 branch_block_stmt_33/merge_stmt_949__exit__
      -- CP-element group 326: 	 branch_block_stmt_33/forx_xend394x_xloopexit_forx_xend394
      -- CP-element group 326: 	 branch_block_stmt_33/if_stmt_943_if_link/$exit
      -- CP-element group 326: 	 branch_block_stmt_33/forx_xbody308_forx_xend394x_xloopexit
      -- CP-element group 326: 	 branch_block_stmt_33/if_stmt_943_if_link/if_choice_transition
      -- CP-element group 326: 	 branch_block_stmt_33/forx_xbody308_forx_xend394x_xloopexit_PhiReq/$entry
      -- CP-element group 326: 	 branch_block_stmt_33/forx_xbody308_forx_xend394x_xloopexit_PhiReq/$exit
      -- CP-element group 326: 	 branch_block_stmt_33/merge_stmt_949_PhiReqMerge
      -- CP-element group 326: 	 branch_block_stmt_33/merge_stmt_949_PhiAck/$entry
      -- CP-element group 326: 	 branch_block_stmt_33/merge_stmt_949_PhiAck/$exit
      -- CP-element group 326: 	 branch_block_stmt_33/merge_stmt_949_PhiAck/dummy
      -- CP-element group 326: 	 branch_block_stmt_33/forx_xend394x_xloopexit_forx_xend394_PhiReq/$entry
      -- CP-element group 326: 	 branch_block_stmt_33/forx_xend394x_xloopexit_forx_xend394_PhiReq/$exit
      -- 
    if_choice_transition_2208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_943_branch_ack_1, ack => convTranspose_CP_39_elements(326)); -- 
    -- CP-element group 327:  fork  transition  place  input  output  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	325 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	523 
    -- CP-element group 327: 	524 
    -- CP-element group 327:  members (12) 
      -- CP-element group 327: 	 branch_block_stmt_33/forx_xbody308_forx_xbody308
      -- CP-element group 327: 	 branch_block_stmt_33/if_stmt_943_else_link/else_choice_transition
      -- CP-element group 327: 	 branch_block_stmt_33/if_stmt_943_else_link/$exit
      -- CP-element group 327: 	 branch_block_stmt_33/forx_xbody308_forx_xbody308_PhiReq/$entry
      -- CP-element group 327: 	 branch_block_stmt_33/forx_xbody308_forx_xbody308_PhiReq/phi_stmt_756/$entry
      -- CP-element group 327: 	 branch_block_stmt_33/forx_xbody308_forx_xbody308_PhiReq/phi_stmt_756/phi_stmt_756_sources/$entry
      -- CP-element group 327: 	 branch_block_stmt_33/forx_xbody308_forx_xbody308_PhiReq/phi_stmt_756/phi_stmt_756_sources/type_cast_762/$entry
      -- CP-element group 327: 	 branch_block_stmt_33/forx_xbody308_forx_xbody308_PhiReq/phi_stmt_756/phi_stmt_756_sources/type_cast_762/SplitProtocol/$entry
      -- CP-element group 327: 	 branch_block_stmt_33/forx_xbody308_forx_xbody308_PhiReq/phi_stmt_756/phi_stmt_756_sources/type_cast_762/SplitProtocol/Sample/$entry
      -- CP-element group 327: 	 branch_block_stmt_33/forx_xbody308_forx_xbody308_PhiReq/phi_stmt_756/phi_stmt_756_sources/type_cast_762/SplitProtocol/Sample/rr
      -- CP-element group 327: 	 branch_block_stmt_33/forx_xbody308_forx_xbody308_PhiReq/phi_stmt_756/phi_stmt_756_sources/type_cast_762/SplitProtocol/Update/$entry
      -- CP-element group 327: 	 branch_block_stmt_33/forx_xbody308_forx_xbody308_PhiReq/phi_stmt_756/phi_stmt_756_sources/type_cast_762/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_943_branch_ack_0, ack => convTranspose_CP_39_elements(327)); -- 
    rr_3714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(327), ack => type_cast_762_inst_req_0); -- 
    cr_3719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(327), ack => type_cast_762_inst_req_1); -- 
    -- CP-element group 328:  transition  input  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	528 
    -- CP-element group 328: successors 
    -- CP-element group 328:  members (3) 
      -- CP-element group 328: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_954_Sample/ra
      -- CP-element group 328: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_954_Sample/$exit
      -- CP-element group 328: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_954_sample_completed_
      -- 
    ra_2226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_954_inst_ack_0, ack => convTranspose_CP_39_elements(328)); -- 
    -- CP-element group 329:  transition  input  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	528 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	334 
    -- CP-element group 329:  members (3) 
      -- CP-element group 329: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_954_Update/ca
      -- CP-element group 329: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_954_Update/$exit
      -- CP-element group 329: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_954_update_completed_
      -- 
    ca_2231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_954_inst_ack_1, ack => convTranspose_CP_39_elements(329)); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	528 
    -- CP-element group 330: successors 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_958_Sample/ra
      -- CP-element group 330: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_958_Sample/$exit
      -- CP-element group 330: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_958_sample_completed_
      -- 
    ra_2240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_958_inst_ack_0, ack => convTranspose_CP_39_elements(330)); -- 
    -- CP-element group 331:  transition  input  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	528 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	334 
    -- CP-element group 331:  members (3) 
      -- CP-element group 331: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_958_Update/$exit
      -- CP-element group 331: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_958_Update/ca
      -- CP-element group 331: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_958_update_completed_
      -- 
    ca_2245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_958_inst_ack_1, ack => convTranspose_CP_39_elements(331)); -- 
    -- CP-element group 332:  transition  input  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	528 
    -- CP-element group 332: successors 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_962_Sample/ra
      -- CP-element group 332: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_962_Sample/$exit
      -- CP-element group 332: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_962_sample_completed_
      -- 
    ra_2254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_962_inst_ack_0, ack => convTranspose_CP_39_elements(332)); -- 
    -- CP-element group 333:  transition  input  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	528 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (3) 
      -- CP-element group 333: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_962_Update/$exit
      -- CP-element group 333: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_962_Update/ca
      -- CP-element group 333: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_962_update_completed_
      -- 
    ca_2259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_962_inst_ack_1, ack => convTranspose_CP_39_elements(333)); -- 
    -- CP-element group 334:  branch  join  transition  place  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	329 
    -- CP-element group 334: 	331 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334: 	336 
    -- CP-element group 334:  members (10) 
      -- CP-element group 334: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979__exit__
      -- CP-element group 334: 	 branch_block_stmt_33/if_stmt_980__entry__
      -- CP-element group 334: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/$exit
      -- CP-element group 334: 	 branch_block_stmt_33/if_stmt_980_else_link/$entry
      -- CP-element group 334: 	 branch_block_stmt_33/if_stmt_980_if_link/$entry
      -- CP-element group 334: 	 branch_block_stmt_33/R_cmp408567_981_place
      -- CP-element group 334: 	 branch_block_stmt_33/if_stmt_980_eval_test/branch_req
      -- CP-element group 334: 	 branch_block_stmt_33/if_stmt_980_eval_test/$exit
      -- CP-element group 334: 	 branch_block_stmt_33/if_stmt_980_eval_test/$entry
      -- CP-element group 334: 	 branch_block_stmt_33/if_stmt_980_dead_link/$entry
      -- 
    branch_req_2267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(334), ack => if_stmt_980_branch_req_0); -- 
    convTranspose_cp_element_group_334: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_334"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(329) & convTranspose_CP_39_elements(331) & convTranspose_CP_39_elements(333);
      gj_convTranspose_cp_element_group_334 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(334), clk => clk, reset => reset); --
    end block;
    -- CP-element group 335:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	337 
    -- CP-element group 335: 	338 
    -- CP-element group 335:  members (18) 
      -- CP-element group 335: 	 branch_block_stmt_33/assign_stmt_992_to_assign_stmt_1021/type_cast_1007_Update/cr
      -- CP-element group 335: 	 branch_block_stmt_33/merge_stmt_986__exit__
      -- CP-element group 335: 	 branch_block_stmt_33/assign_stmt_992_to_assign_stmt_1021__entry__
      -- CP-element group 335: 	 branch_block_stmt_33/assign_stmt_992_to_assign_stmt_1021/type_cast_1007_sample_start_
      -- CP-element group 335: 	 branch_block_stmt_33/assign_stmt_992_to_assign_stmt_1021/$entry
      -- CP-element group 335: 	 branch_block_stmt_33/assign_stmt_992_to_assign_stmt_1021/type_cast_1007_update_start_
      -- CP-element group 335: 	 branch_block_stmt_33/assign_stmt_992_to_assign_stmt_1021/type_cast_1007_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_33/forx_xend394_bbx_xnph569
      -- CP-element group 335: 	 branch_block_stmt_33/if_stmt_980_if_link/if_choice_transition
      -- CP-element group 335: 	 branch_block_stmt_33/assign_stmt_992_to_assign_stmt_1021/type_cast_1007_Sample/rr
      -- CP-element group 335: 	 branch_block_stmt_33/if_stmt_980_if_link/$exit
      -- CP-element group 335: 	 branch_block_stmt_33/assign_stmt_992_to_assign_stmt_1021/type_cast_1007_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_33/forx_xend394_bbx_xnph569_PhiReq/$entry
      -- CP-element group 335: 	 branch_block_stmt_33/forx_xend394_bbx_xnph569_PhiReq/$exit
      -- CP-element group 335: 	 branch_block_stmt_33/merge_stmt_986_PhiReqMerge
      -- CP-element group 335: 	 branch_block_stmt_33/merge_stmt_986_PhiAck/$entry
      -- CP-element group 335: 	 branch_block_stmt_33/merge_stmt_986_PhiAck/$exit
      -- CP-element group 335: 	 branch_block_stmt_33/merge_stmt_986_PhiAck/dummy
      -- 
    if_choice_transition_2272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_980_branch_ack_1, ack => convTranspose_CP_39_elements(335)); -- 
    cr_2294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(335), ack => type_cast_1007_inst_req_1); -- 
    rr_2289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(335), ack => type_cast_1007_inst_req_0); -- 
    -- CP-element group 336:  transition  place  input  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	334 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	535 
    -- CP-element group 336:  members (5) 
      -- CP-element group 336: 	 branch_block_stmt_33/forx_xend394_forx_xend417
      -- CP-element group 336: 	 branch_block_stmt_33/if_stmt_980_else_link/else_choice_transition
      -- CP-element group 336: 	 branch_block_stmt_33/if_stmt_980_else_link/$exit
      -- CP-element group 336: 	 branch_block_stmt_33/forx_xend394_forx_xend417_PhiReq/$entry
      -- CP-element group 336: 	 branch_block_stmt_33/forx_xend394_forx_xend417_PhiReq/$exit
      -- 
    else_choice_transition_2276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_980_branch_ack_0, ack => convTranspose_CP_39_elements(336)); -- 
    -- CP-element group 337:  transition  input  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	335 
    -- CP-element group 337: successors 
    -- CP-element group 337:  members (3) 
      -- CP-element group 337: 	 branch_block_stmt_33/assign_stmt_992_to_assign_stmt_1021/type_cast_1007_sample_completed_
      -- CP-element group 337: 	 branch_block_stmt_33/assign_stmt_992_to_assign_stmt_1021/type_cast_1007_Sample/ra
      -- CP-element group 337: 	 branch_block_stmt_33/assign_stmt_992_to_assign_stmt_1021/type_cast_1007_Sample/$exit
      -- 
    ra_2290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1007_inst_ack_0, ack => convTranspose_CP_39_elements(337)); -- 
    -- CP-element group 338:  transition  place  input  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	335 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	529 
    -- CP-element group 338:  members (9) 
      -- CP-element group 338: 	 branch_block_stmt_33/assign_stmt_992_to_assign_stmt_1021/type_cast_1007_Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_33/assign_stmt_992_to_assign_stmt_1021__exit__
      -- CP-element group 338: 	 branch_block_stmt_33/bbx_xnph569_forx_xbody410
      -- CP-element group 338: 	 branch_block_stmt_33/assign_stmt_992_to_assign_stmt_1021/type_cast_1007_Update/ca
      -- CP-element group 338: 	 branch_block_stmt_33/assign_stmt_992_to_assign_stmt_1021/$exit
      -- CP-element group 338: 	 branch_block_stmt_33/assign_stmt_992_to_assign_stmt_1021/type_cast_1007_update_completed_
      -- CP-element group 338: 	 branch_block_stmt_33/bbx_xnph569_forx_xbody410_PhiReq/$entry
      -- CP-element group 338: 	 branch_block_stmt_33/bbx_xnph569_forx_xbody410_PhiReq/phi_stmt_1024/$entry
      -- CP-element group 338: 	 branch_block_stmt_33/bbx_xnph569_forx_xbody410_PhiReq/phi_stmt_1024/phi_stmt_1024_sources/$entry
      -- 
    ca_2295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1007_inst_ack_1, ack => convTranspose_CP_39_elements(338)); -- 
    -- CP-element group 339:  transition  input  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	534 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	345 
    -- CP-element group 339:  members (3) 
      -- CP-element group 339: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_final_index_sum_regn_Sample/ack
      -- CP-element group 339: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_final_index_sum_regn_Sample/$exit
      -- CP-element group 339: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_final_index_sum_regn_sample_complete
      -- 
    ack_2324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1036_index_offset_ack_0, ack => convTranspose_CP_39_elements(339)); -- 
    -- CP-element group 340:  transition  input  output  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	534 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (11) 
      -- CP-element group 340: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_final_index_sum_regn_Update/$exit
      -- CP-element group 340: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/addr_of_1037_request/req
      -- CP-element group 340: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_base_plus_offset/sum_rename_req
      -- CP-element group 340: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_final_index_sum_regn_Update/ack
      -- CP-element group 340: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_base_plus_offset/$exit
      -- CP-element group 340: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/addr_of_1037_request/$entry
      -- CP-element group 340: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_base_plus_offset/$entry
      -- CP-element group 340: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_offset_calculated
      -- CP-element group 340: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_root_address_calculated
      -- CP-element group 340: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/addr_of_1037_sample_start_
      -- CP-element group 340: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_base_plus_offset/sum_rename_ack
      -- 
    ack_2329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1036_index_offset_ack_1, ack => convTranspose_CP_39_elements(340)); -- 
    req_2338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(340), ack => addr_of_1037_final_reg_req_0); -- 
    -- CP-element group 341:  transition  input  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341:  members (3) 
      -- CP-element group 341: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/addr_of_1037_request/$exit
      -- CP-element group 341: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/addr_of_1037_request/ack
      -- CP-element group 341: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/addr_of_1037_sample_completed_
      -- 
    ack_2339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1037_final_reg_ack_0, ack => convTranspose_CP_39_elements(341)); -- 
    -- CP-element group 342:  join  fork  transition  input  output  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	534 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	343 
    -- CP-element group 342:  members (28) 
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_base_addr_resize/$exit
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_sample_start_
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_base_address_resized
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_root_address_calculated
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_word_address_calculated
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_base_address_calculated
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/addr_of_1037_complete/ack
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/addr_of_1037_complete/$exit
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/addr_of_1037_update_completed_
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_base_addr_resize/$entry
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_base_addr_resize/base_resize_req
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_base_addr_resize/base_resize_ack
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_base_plus_offset/$entry
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_base_plus_offset/$exit
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_base_plus_offset/sum_rename_req
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_base_plus_offset/sum_rename_ack
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_word_addrgen/$entry
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_word_addrgen/$exit
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_word_addrgen/root_register_req
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_word_addrgen/root_register_ack
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_Sample/ptr_deref_1040_Split/$entry
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_Sample/ptr_deref_1040_Split/$exit
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_Sample/ptr_deref_1040_Split/split_req
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_Sample/ptr_deref_1040_Split/split_ack
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_Sample/word_access_start/$entry
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_Sample/word_access_start/word_0/$entry
      -- CP-element group 342: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_Sample/word_access_start/word_0/rr
      -- 
    ack_2344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1037_final_reg_ack_1, ack => convTranspose_CP_39_elements(342)); -- 
    rr_2382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(342), ack => ptr_deref_1040_store_0_req_0); -- 
    -- CP-element group 343:  transition  input  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	342 
    -- CP-element group 343: successors 
    -- CP-element group 343:  members (5) 
      -- CP-element group 343: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_sample_completed_
      -- CP-element group 343: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_Sample/$exit
      -- CP-element group 343: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_Sample/word_access_start/$exit
      -- CP-element group 343: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_Sample/word_access_start/word_0/$exit
      -- CP-element group 343: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_Sample/word_access_start/word_0/ra
      -- 
    ra_2383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1040_store_0_ack_0, ack => convTranspose_CP_39_elements(343)); -- 
    -- CP-element group 344:  transition  input  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	534 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	345 
    -- CP-element group 344:  members (5) 
      -- CP-element group 344: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_Update/$exit
      -- CP-element group 344: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_Update/word_access_complete/$exit
      -- CP-element group 344: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_Update/word_access_complete/word_0/$exit
      -- CP-element group 344: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_Update/word_access_complete/word_0/ca
      -- 
    ca_2394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1040_store_0_ack_1, ack => convTranspose_CP_39_elements(344)); -- 
    -- CP-element group 345:  branch  join  transition  place  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	339 
    -- CP-element group 345: 	344 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345: 	347 
    -- CP-element group 345:  members (10) 
      -- CP-element group 345: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054__exit__
      -- CP-element group 345: 	 branch_block_stmt_33/if_stmt_1055__entry__
      -- CP-element group 345: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/$exit
      -- CP-element group 345: 	 branch_block_stmt_33/if_stmt_1055_dead_link/$entry
      -- CP-element group 345: 	 branch_block_stmt_33/if_stmt_1055_eval_test/$entry
      -- CP-element group 345: 	 branch_block_stmt_33/if_stmt_1055_eval_test/$exit
      -- CP-element group 345: 	 branch_block_stmt_33/if_stmt_1055_eval_test/branch_req
      -- CP-element group 345: 	 branch_block_stmt_33/R_exitcond_1056_place
      -- CP-element group 345: 	 branch_block_stmt_33/if_stmt_1055_if_link/$entry
      -- CP-element group 345: 	 branch_block_stmt_33/if_stmt_1055_else_link/$entry
      -- 
    branch_req_2402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(345), ack => if_stmt_1055_branch_req_0); -- 
    convTranspose_cp_element_group_345: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_345"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(339) & convTranspose_CP_39_elements(344);
      gj_convTranspose_cp_element_group_345 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(345), clk => clk, reset => reset); --
    end block;
    -- CP-element group 346:  merge  transition  place  input  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	535 
    -- CP-element group 346:  members (13) 
      -- CP-element group 346: 	 branch_block_stmt_33/merge_stmt_1061__exit__
      -- CP-element group 346: 	 branch_block_stmt_33/forx_xend417x_xloopexit_forx_xend417
      -- CP-element group 346: 	 branch_block_stmt_33/if_stmt_1055_if_link/$exit
      -- CP-element group 346: 	 branch_block_stmt_33/if_stmt_1055_if_link/if_choice_transition
      -- CP-element group 346: 	 branch_block_stmt_33/forx_xbody410_forx_xend417x_xloopexit
      -- CP-element group 346: 	 branch_block_stmt_33/forx_xbody410_forx_xend417x_xloopexit_PhiReq/$entry
      -- CP-element group 346: 	 branch_block_stmt_33/forx_xbody410_forx_xend417x_xloopexit_PhiReq/$exit
      -- CP-element group 346: 	 branch_block_stmt_33/merge_stmt_1061_PhiReqMerge
      -- CP-element group 346: 	 branch_block_stmt_33/merge_stmt_1061_PhiAck/$entry
      -- CP-element group 346: 	 branch_block_stmt_33/merge_stmt_1061_PhiAck/$exit
      -- CP-element group 346: 	 branch_block_stmt_33/merge_stmt_1061_PhiAck/dummy
      -- CP-element group 346: 	 branch_block_stmt_33/forx_xend417x_xloopexit_forx_xend417_PhiReq/$entry
      -- CP-element group 346: 	 branch_block_stmt_33/forx_xend417x_xloopexit_forx_xend417_PhiReq/$exit
      -- 
    if_choice_transition_2407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1055_branch_ack_1, ack => convTranspose_CP_39_elements(346)); -- 
    -- CP-element group 347:  fork  transition  place  input  output  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	345 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	530 
    -- CP-element group 347: 	531 
    -- CP-element group 347:  members (12) 
      -- CP-element group 347: 	 branch_block_stmt_33/if_stmt_1055_else_link/$exit
      -- CP-element group 347: 	 branch_block_stmt_33/if_stmt_1055_else_link/else_choice_transition
      -- CP-element group 347: 	 branch_block_stmt_33/forx_xbody410_forx_xbody410
      -- CP-element group 347: 	 branch_block_stmt_33/forx_xbody410_forx_xbody410_PhiReq/$entry
      -- CP-element group 347: 	 branch_block_stmt_33/forx_xbody410_forx_xbody410_PhiReq/phi_stmt_1024/$entry
      -- CP-element group 347: 	 branch_block_stmt_33/forx_xbody410_forx_xbody410_PhiReq/phi_stmt_1024/phi_stmt_1024_sources/$entry
      -- CP-element group 347: 	 branch_block_stmt_33/forx_xbody410_forx_xbody410_PhiReq/phi_stmt_1024/phi_stmt_1024_sources/type_cast_1030/$entry
      -- CP-element group 347: 	 branch_block_stmt_33/forx_xbody410_forx_xbody410_PhiReq/phi_stmt_1024/phi_stmt_1024_sources/type_cast_1030/SplitProtocol/$entry
      -- CP-element group 347: 	 branch_block_stmt_33/forx_xbody410_forx_xbody410_PhiReq/phi_stmt_1024/phi_stmt_1024_sources/type_cast_1030/SplitProtocol/Sample/$entry
      -- CP-element group 347: 	 branch_block_stmt_33/forx_xbody410_forx_xbody410_PhiReq/phi_stmt_1024/phi_stmt_1024_sources/type_cast_1030/SplitProtocol/Sample/rr
      -- CP-element group 347: 	 branch_block_stmt_33/forx_xbody410_forx_xbody410_PhiReq/phi_stmt_1024/phi_stmt_1024_sources/type_cast_1030/SplitProtocol/Update/$entry
      -- CP-element group 347: 	 branch_block_stmt_33/forx_xbody410_forx_xbody410_PhiReq/phi_stmt_1024/phi_stmt_1024_sources/type_cast_1030/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1055_branch_ack_0, ack => convTranspose_CP_39_elements(347)); -- 
    rr_3791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(347), ack => type_cast_1030_inst_req_0); -- 
    cr_3796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(347), ack => type_cast_1030_inst_req_1); -- 
    -- CP-element group 348:  transition  input  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	535 
    -- CP-element group 348: successors 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/call_stmt_1066_sample_completed_
      -- CP-element group 348: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/call_stmt_1066_Sample/$exit
      -- CP-element group 348: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/call_stmt_1066_Sample/cra
      -- 
    cra_2425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1066_call_ack_0, ack => convTranspose_CP_39_elements(348)); -- 
    -- CP-element group 349:  transition  input  output  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	535 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	350 
    -- CP-element group 349:  members (6) 
      -- CP-element group 349: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/call_stmt_1066_update_completed_
      -- CP-element group 349: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/call_stmt_1066_Update/$exit
      -- CP-element group 349: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/call_stmt_1066_Update/cca
      -- CP-element group 349: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/type_cast_1071_sample_start_
      -- CP-element group 349: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/type_cast_1071_Sample/$entry
      -- CP-element group 349: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/type_cast_1071_Sample/rr
      -- 
    cca_2430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1066_call_ack_1, ack => convTranspose_CP_39_elements(349)); -- 
    rr_2438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(349), ack => type_cast_1071_inst_req_0); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	349 
    -- CP-element group 350: successors 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/type_cast_1071_sample_completed_
      -- CP-element group 350: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/type_cast_1071_Sample/$exit
      -- CP-element group 350: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/type_cast_1071_Sample/ra
      -- 
    ra_2439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1071_inst_ack_0, ack => convTranspose_CP_39_elements(350)); -- 
    -- CP-element group 351:  transition  input  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	535 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	456 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/type_cast_1071_update_completed_
      -- CP-element group 351: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/type_cast_1071_Update/$exit
      -- CP-element group 351: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/type_cast_1071_Update/ca
      -- 
    ca_2444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1071_inst_ack_1, ack => convTranspose_CP_39_elements(351)); -- 
    -- CP-element group 352:  transition  input  output  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	535 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (6) 
      -- CP-element group 352: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1073_sample_completed_
      -- CP-element group 352: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1073_update_start_
      -- CP-element group 352: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1073_Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1073_Sample/ack
      -- CP-element group 352: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1073_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1073_Update/req
      -- 
    ack_2453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1073_inst_ack_0, ack => convTranspose_CP_39_elements(352)); -- 
    req_2457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(352), ack => WPIPE_Block0_start_1073_inst_req_1); -- 
    -- CP-element group 353:  transition  input  output  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	354 
    -- CP-element group 353:  members (6) 
      -- CP-element group 353: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1073_update_completed_
      -- CP-element group 353: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1073_Update/$exit
      -- CP-element group 353: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1073_Update/ack
      -- CP-element group 353: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1076_sample_start_
      -- CP-element group 353: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1076_Sample/$entry
      -- CP-element group 353: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1076_Sample/req
      -- 
    ack_2458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1073_inst_ack_1, ack => convTranspose_CP_39_elements(353)); -- 
    req_2466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(353), ack => WPIPE_Block0_start_1076_inst_req_0); -- 
    -- CP-element group 354:  transition  input  output  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	353 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	355 
    -- CP-element group 354:  members (6) 
      -- CP-element group 354: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1076_sample_completed_
      -- CP-element group 354: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1076_update_start_
      -- CP-element group 354: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1076_Sample/$exit
      -- CP-element group 354: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1076_Sample/ack
      -- CP-element group 354: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1076_Update/$entry
      -- CP-element group 354: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1076_Update/req
      -- 
    ack_2467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1076_inst_ack_0, ack => convTranspose_CP_39_elements(354)); -- 
    req_2471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(354), ack => WPIPE_Block0_start_1076_inst_req_1); -- 
    -- CP-element group 355:  transition  input  output  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	354 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (6) 
      -- CP-element group 355: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1076_update_completed_
      -- CP-element group 355: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1076_Update/$exit
      -- CP-element group 355: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1076_Update/ack
      -- CP-element group 355: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1079_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1079_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1079_Sample/req
      -- 
    ack_2472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1076_inst_ack_1, ack => convTranspose_CP_39_elements(355)); -- 
    req_2480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(355), ack => WPIPE_Block0_start_1079_inst_req_0); -- 
    -- CP-element group 356:  transition  input  output  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	357 
    -- CP-element group 356:  members (6) 
      -- CP-element group 356: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1079_sample_completed_
      -- CP-element group 356: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1079_update_start_
      -- CP-element group 356: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1079_Sample/$exit
      -- CP-element group 356: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1079_Sample/ack
      -- CP-element group 356: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1079_Update/$entry
      -- CP-element group 356: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1079_Update/req
      -- 
    ack_2481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1079_inst_ack_0, ack => convTranspose_CP_39_elements(356)); -- 
    req_2485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(356), ack => WPIPE_Block0_start_1079_inst_req_1); -- 
    -- CP-element group 357:  transition  input  output  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	356 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (6) 
      -- CP-element group 357: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1079_update_completed_
      -- CP-element group 357: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1079_Update/$exit
      -- CP-element group 357: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1079_Update/ack
      -- CP-element group 357: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1082_sample_start_
      -- CP-element group 357: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1082_Sample/$entry
      -- CP-element group 357: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1082_Sample/req
      -- 
    ack_2486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1079_inst_ack_1, ack => convTranspose_CP_39_elements(357)); -- 
    req_2494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(357), ack => WPIPE_Block0_start_1082_inst_req_0); -- 
    -- CP-element group 358:  transition  input  output  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (6) 
      -- CP-element group 358: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1082_sample_completed_
      -- CP-element group 358: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1082_update_start_
      -- CP-element group 358: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1082_Sample/$exit
      -- CP-element group 358: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1082_Sample/ack
      -- CP-element group 358: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1082_Update/$entry
      -- CP-element group 358: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1082_Update/req
      -- 
    ack_2495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1082_inst_ack_0, ack => convTranspose_CP_39_elements(358)); -- 
    req_2499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(358), ack => WPIPE_Block0_start_1082_inst_req_1); -- 
    -- CP-element group 359:  transition  input  output  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	360 
    -- CP-element group 359:  members (6) 
      -- CP-element group 359: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1082_update_completed_
      -- CP-element group 359: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1082_Update/$exit
      -- CP-element group 359: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1082_Update/ack
      -- CP-element group 359: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1085_sample_start_
      -- CP-element group 359: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1085_Sample/$entry
      -- CP-element group 359: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1085_Sample/req
      -- 
    ack_2500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1082_inst_ack_1, ack => convTranspose_CP_39_elements(359)); -- 
    req_2508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(359), ack => WPIPE_Block0_start_1085_inst_req_0); -- 
    -- CP-element group 360:  transition  input  output  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	359 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360:  members (6) 
      -- CP-element group 360: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1085_sample_completed_
      -- CP-element group 360: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1085_update_start_
      -- CP-element group 360: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1085_Sample/$exit
      -- CP-element group 360: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1085_Sample/ack
      -- CP-element group 360: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1085_Update/$entry
      -- CP-element group 360: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1085_Update/req
      -- 
    ack_2509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1085_inst_ack_0, ack => convTranspose_CP_39_elements(360)); -- 
    req_2513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(360), ack => WPIPE_Block0_start_1085_inst_req_1); -- 
    -- CP-element group 361:  transition  input  output  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	360 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (6) 
      -- CP-element group 361: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1085_update_completed_
      -- CP-element group 361: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1085_Update/$exit
      -- CP-element group 361: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1085_Update/ack
      -- CP-element group 361: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1088_sample_start_
      -- CP-element group 361: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1088_Sample/$entry
      -- CP-element group 361: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1088_Sample/req
      -- 
    ack_2514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1085_inst_ack_1, ack => convTranspose_CP_39_elements(361)); -- 
    req_2522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(361), ack => WPIPE_Block0_start_1088_inst_req_0); -- 
    -- CP-element group 362:  transition  input  output  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362:  members (6) 
      -- CP-element group 362: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1088_sample_completed_
      -- CP-element group 362: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1088_update_start_
      -- CP-element group 362: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1088_Sample/$exit
      -- CP-element group 362: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1088_Sample/ack
      -- CP-element group 362: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1088_Update/$entry
      -- CP-element group 362: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1088_Update/req
      -- 
    ack_2523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1088_inst_ack_0, ack => convTranspose_CP_39_elements(362)); -- 
    req_2527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(362), ack => WPIPE_Block0_start_1088_inst_req_1); -- 
    -- CP-element group 363:  transition  input  output  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (6) 
      -- CP-element group 363: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1088_update_completed_
      -- CP-element group 363: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1088_Update/$exit
      -- CP-element group 363: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1088_Update/ack
      -- CP-element group 363: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1091_sample_start_
      -- CP-element group 363: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1091_Sample/$entry
      -- CP-element group 363: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1091_Sample/req
      -- 
    ack_2528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1088_inst_ack_1, ack => convTranspose_CP_39_elements(363)); -- 
    req_2536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(363), ack => WPIPE_Block0_start_1091_inst_req_0); -- 
    -- CP-element group 364:  transition  input  output  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	365 
    -- CP-element group 364:  members (6) 
      -- CP-element group 364: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1091_sample_completed_
      -- CP-element group 364: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1091_update_start_
      -- CP-element group 364: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1091_Sample/$exit
      -- CP-element group 364: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1091_Sample/ack
      -- CP-element group 364: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1091_Update/$entry
      -- CP-element group 364: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1091_Update/req
      -- 
    ack_2537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1091_inst_ack_0, ack => convTranspose_CP_39_elements(364)); -- 
    req_2541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(364), ack => WPIPE_Block0_start_1091_inst_req_1); -- 
    -- CP-element group 365:  transition  input  output  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	364 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365:  members (6) 
      -- CP-element group 365: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1091_update_completed_
      -- CP-element group 365: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1091_Update/$exit
      -- CP-element group 365: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1091_Update/ack
      -- CP-element group 365: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1094_sample_start_
      -- CP-element group 365: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1094_Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1094_Sample/req
      -- 
    ack_2542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1091_inst_ack_1, ack => convTranspose_CP_39_elements(365)); -- 
    req_2550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(365), ack => WPIPE_Block0_start_1094_inst_req_0); -- 
    -- CP-element group 366:  transition  input  output  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	367 
    -- CP-element group 366:  members (6) 
      -- CP-element group 366: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1094_sample_completed_
      -- CP-element group 366: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1094_update_start_
      -- CP-element group 366: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1094_Sample/$exit
      -- CP-element group 366: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1094_Sample/ack
      -- CP-element group 366: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1094_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1094_Update/req
      -- 
    ack_2551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1094_inst_ack_0, ack => convTranspose_CP_39_elements(366)); -- 
    req_2555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(366), ack => WPIPE_Block0_start_1094_inst_req_1); -- 
    -- CP-element group 367:  transition  input  output  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	366 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367:  members (6) 
      -- CP-element group 367: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1094_update_completed_
      -- CP-element group 367: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1094_Update/$exit
      -- CP-element group 367: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1094_Update/ack
      -- CP-element group 367: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1097_sample_start_
      -- CP-element group 367: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1097_Sample/$entry
      -- CP-element group 367: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1097_Sample/req
      -- 
    ack_2556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1094_inst_ack_1, ack => convTranspose_CP_39_elements(367)); -- 
    req_2564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(367), ack => WPIPE_Block0_start_1097_inst_req_0); -- 
    -- CP-element group 368:  transition  input  output  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	369 
    -- CP-element group 368:  members (6) 
      -- CP-element group 368: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1097_sample_completed_
      -- CP-element group 368: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1097_update_start_
      -- CP-element group 368: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1097_Sample/$exit
      -- CP-element group 368: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1097_Sample/ack
      -- CP-element group 368: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1097_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1097_Update/req
      -- 
    ack_2565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1097_inst_ack_0, ack => convTranspose_CP_39_elements(368)); -- 
    req_2569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(368), ack => WPIPE_Block0_start_1097_inst_req_1); -- 
    -- CP-element group 369:  transition  input  output  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	368 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	370 
    -- CP-element group 369:  members (6) 
      -- CP-element group 369: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1097_update_completed_
      -- CP-element group 369: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1097_Update/$exit
      -- CP-element group 369: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1097_Update/ack
      -- CP-element group 369: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1100_sample_start_
      -- CP-element group 369: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1100_Sample/$entry
      -- CP-element group 369: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1100_Sample/req
      -- 
    ack_2570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1097_inst_ack_1, ack => convTranspose_CP_39_elements(369)); -- 
    req_2578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(369), ack => WPIPE_Block0_start_1100_inst_req_0); -- 
    -- CP-element group 370:  transition  input  output  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	369 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	371 
    -- CP-element group 370:  members (6) 
      -- CP-element group 370: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1100_sample_completed_
      -- CP-element group 370: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1100_update_start_
      -- CP-element group 370: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1100_Sample/$exit
      -- CP-element group 370: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1100_Sample/ack
      -- CP-element group 370: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1100_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1100_Update/req
      -- 
    ack_2579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1100_inst_ack_0, ack => convTranspose_CP_39_elements(370)); -- 
    req_2583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(370), ack => WPIPE_Block0_start_1100_inst_req_1); -- 
    -- CP-element group 371:  transition  input  output  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	370 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (6) 
      -- CP-element group 371: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1100_update_completed_
      -- CP-element group 371: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1100_Update/$exit
      -- CP-element group 371: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1100_Update/ack
      -- CP-element group 371: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1103_sample_start_
      -- CP-element group 371: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1103_Sample/$entry
      -- CP-element group 371: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1103_Sample/req
      -- 
    ack_2584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1100_inst_ack_1, ack => convTranspose_CP_39_elements(371)); -- 
    req_2592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(371), ack => WPIPE_Block0_start_1103_inst_req_0); -- 
    -- CP-element group 372:  transition  input  output  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (6) 
      -- CP-element group 372: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1103_sample_completed_
      -- CP-element group 372: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1103_update_start_
      -- CP-element group 372: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1103_Sample/$exit
      -- CP-element group 372: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1103_Sample/ack
      -- CP-element group 372: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1103_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1103_Update/req
      -- 
    ack_2593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1103_inst_ack_0, ack => convTranspose_CP_39_elements(372)); -- 
    req_2597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(372), ack => WPIPE_Block0_start_1103_inst_req_1); -- 
    -- CP-element group 373:  transition  input  output  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (6) 
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1103_update_completed_
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1103_Update/$exit
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1103_Update/ack
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1106_sample_start_
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1106_Sample/$entry
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1106_Sample/req
      -- 
    ack_2598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1103_inst_ack_1, ack => convTranspose_CP_39_elements(373)); -- 
    req_2606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => WPIPE_Block0_start_1106_inst_req_0); -- 
    -- CP-element group 374:  transition  input  output  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	375 
    -- CP-element group 374:  members (6) 
      -- CP-element group 374: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1106_sample_completed_
      -- CP-element group 374: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1106_update_start_
      -- CP-element group 374: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1106_Sample/$exit
      -- CP-element group 374: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1106_Sample/ack
      -- CP-element group 374: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1106_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1106_Update/req
      -- 
    ack_2607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1106_inst_ack_0, ack => convTranspose_CP_39_elements(374)); -- 
    req_2611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(374), ack => WPIPE_Block0_start_1106_inst_req_1); -- 
    -- CP-element group 375:  transition  input  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	374 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	456 
    -- CP-element group 375:  members (3) 
      -- CP-element group 375: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1106_update_completed_
      -- CP-element group 375: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1106_Update/$exit
      -- CP-element group 375: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1106_Update/ack
      -- 
    ack_2612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1106_inst_ack_1, ack => convTranspose_CP_39_elements(375)); -- 
    -- CP-element group 376:  transition  input  output  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	535 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	377 
    -- CP-element group 376:  members (6) 
      -- CP-element group 376: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1109_sample_completed_
      -- CP-element group 376: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1109_update_start_
      -- CP-element group 376: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1109_Sample/$exit
      -- CP-element group 376: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1109_Sample/ack
      -- CP-element group 376: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1109_Update/$entry
      -- CP-element group 376: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1109_Update/req
      -- 
    ack_2621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1109_inst_ack_0, ack => convTranspose_CP_39_elements(376)); -- 
    req_2625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(376), ack => WPIPE_Block1_start_1109_inst_req_1); -- 
    -- CP-element group 377:  transition  input  output  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	376 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	378 
    -- CP-element group 377:  members (6) 
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1109_update_completed_
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1109_Update/$exit
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1109_Update/ack
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1112_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1112_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1112_Sample/req
      -- 
    ack_2626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1109_inst_ack_1, ack => convTranspose_CP_39_elements(377)); -- 
    req_2634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => WPIPE_Block1_start_1112_inst_req_0); -- 
    -- CP-element group 378:  transition  input  output  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	377 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	379 
    -- CP-element group 378:  members (6) 
      -- CP-element group 378: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1112_sample_completed_
      -- CP-element group 378: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1112_update_start_
      -- CP-element group 378: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1112_Sample/$exit
      -- CP-element group 378: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1112_Sample/ack
      -- CP-element group 378: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1112_Update/$entry
      -- CP-element group 378: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1112_Update/req
      -- 
    ack_2635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1112_inst_ack_0, ack => convTranspose_CP_39_elements(378)); -- 
    req_2639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(378), ack => WPIPE_Block1_start_1112_inst_req_1); -- 
    -- CP-element group 379:  transition  input  output  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	378 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	380 
    -- CP-element group 379:  members (6) 
      -- CP-element group 379: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1112_update_completed_
      -- CP-element group 379: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1112_Update/$exit
      -- CP-element group 379: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1112_Update/ack
      -- CP-element group 379: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1115_sample_start_
      -- CP-element group 379: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1115_Sample/$entry
      -- CP-element group 379: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1115_Sample/req
      -- 
    ack_2640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1112_inst_ack_1, ack => convTranspose_CP_39_elements(379)); -- 
    req_2648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(379), ack => WPIPE_Block1_start_1115_inst_req_0); -- 
    -- CP-element group 380:  transition  input  output  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	379 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	381 
    -- CP-element group 380:  members (6) 
      -- CP-element group 380: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1115_sample_completed_
      -- CP-element group 380: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1115_update_start_
      -- CP-element group 380: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1115_Sample/$exit
      -- CP-element group 380: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1115_Sample/ack
      -- CP-element group 380: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1115_Update/$entry
      -- CP-element group 380: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1115_Update/req
      -- 
    ack_2649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1115_inst_ack_0, ack => convTranspose_CP_39_elements(380)); -- 
    req_2653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(380), ack => WPIPE_Block1_start_1115_inst_req_1); -- 
    -- CP-element group 381:  transition  input  output  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	380 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	382 
    -- CP-element group 381:  members (6) 
      -- CP-element group 381: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1115_update_completed_
      -- CP-element group 381: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1115_Update/$exit
      -- CP-element group 381: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1115_Update/ack
      -- CP-element group 381: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1118_sample_start_
      -- CP-element group 381: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1118_Sample/$entry
      -- CP-element group 381: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1118_Sample/req
      -- 
    ack_2654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1115_inst_ack_1, ack => convTranspose_CP_39_elements(381)); -- 
    req_2662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(381), ack => WPIPE_Block1_start_1118_inst_req_0); -- 
    -- CP-element group 382:  transition  input  output  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	381 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	383 
    -- CP-element group 382:  members (6) 
      -- CP-element group 382: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1118_sample_completed_
      -- CP-element group 382: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1118_update_start_
      -- CP-element group 382: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1118_Sample/$exit
      -- CP-element group 382: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1118_Sample/ack
      -- CP-element group 382: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1118_Update/$entry
      -- CP-element group 382: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1118_Update/req
      -- 
    ack_2663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1118_inst_ack_0, ack => convTranspose_CP_39_elements(382)); -- 
    req_2667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(382), ack => WPIPE_Block1_start_1118_inst_req_1); -- 
    -- CP-element group 383:  transition  input  output  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	382 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	384 
    -- CP-element group 383:  members (6) 
      -- CP-element group 383: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1118_update_completed_
      -- CP-element group 383: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1118_Update/$exit
      -- CP-element group 383: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1118_Update/ack
      -- CP-element group 383: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1121_sample_start_
      -- CP-element group 383: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1121_Sample/$entry
      -- CP-element group 383: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1121_Sample/req
      -- 
    ack_2668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1118_inst_ack_1, ack => convTranspose_CP_39_elements(383)); -- 
    req_2676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(383), ack => WPIPE_Block1_start_1121_inst_req_0); -- 
    -- CP-element group 384:  transition  input  output  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	383 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	385 
    -- CP-element group 384:  members (6) 
      -- CP-element group 384: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1121_sample_completed_
      -- CP-element group 384: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1121_update_start_
      -- CP-element group 384: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1121_Sample/$exit
      -- CP-element group 384: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1121_Sample/ack
      -- CP-element group 384: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1121_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1121_Update/req
      -- 
    ack_2677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1121_inst_ack_0, ack => convTranspose_CP_39_elements(384)); -- 
    req_2681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(384), ack => WPIPE_Block1_start_1121_inst_req_1); -- 
    -- CP-element group 385:  transition  input  output  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	384 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	386 
    -- CP-element group 385:  members (6) 
      -- CP-element group 385: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1121_update_completed_
      -- CP-element group 385: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1121_Update/$exit
      -- CP-element group 385: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1121_Update/ack
      -- CP-element group 385: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1124_sample_start_
      -- CP-element group 385: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1124_Sample/$entry
      -- CP-element group 385: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1124_Sample/req
      -- 
    ack_2682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1121_inst_ack_1, ack => convTranspose_CP_39_elements(385)); -- 
    req_2690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(385), ack => WPIPE_Block1_start_1124_inst_req_0); -- 
    -- CP-element group 386:  transition  input  output  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	385 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	387 
    -- CP-element group 386:  members (6) 
      -- CP-element group 386: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1124_sample_completed_
      -- CP-element group 386: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1124_update_start_
      -- CP-element group 386: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1124_Sample/$exit
      -- CP-element group 386: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1124_Sample/ack
      -- CP-element group 386: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1124_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1124_Update/req
      -- 
    ack_2691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1124_inst_ack_0, ack => convTranspose_CP_39_elements(386)); -- 
    req_2695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(386), ack => WPIPE_Block1_start_1124_inst_req_1); -- 
    -- CP-element group 387:  transition  input  output  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	386 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	388 
    -- CP-element group 387:  members (6) 
      -- CP-element group 387: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1124_update_completed_
      -- CP-element group 387: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1124_Update/$exit
      -- CP-element group 387: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1124_Update/ack
      -- CP-element group 387: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1127_sample_start_
      -- CP-element group 387: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1127_Sample/$entry
      -- CP-element group 387: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1127_Sample/req
      -- 
    ack_2696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1124_inst_ack_1, ack => convTranspose_CP_39_elements(387)); -- 
    req_2704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(387), ack => WPIPE_Block1_start_1127_inst_req_0); -- 
    -- CP-element group 388:  transition  input  output  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	387 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	389 
    -- CP-element group 388:  members (6) 
      -- CP-element group 388: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1127_sample_completed_
      -- CP-element group 388: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1127_update_start_
      -- CP-element group 388: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1127_Sample/$exit
      -- CP-element group 388: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1127_Sample/ack
      -- CP-element group 388: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1127_Update/$entry
      -- CP-element group 388: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1127_Update/req
      -- 
    ack_2705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1127_inst_ack_0, ack => convTranspose_CP_39_elements(388)); -- 
    req_2709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(388), ack => WPIPE_Block1_start_1127_inst_req_1); -- 
    -- CP-element group 389:  transition  input  output  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	388 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	390 
    -- CP-element group 389:  members (6) 
      -- CP-element group 389: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1127_update_completed_
      -- CP-element group 389: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1127_Update/$exit
      -- CP-element group 389: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1127_Update/ack
      -- CP-element group 389: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1130_sample_start_
      -- CP-element group 389: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1130_Sample/$entry
      -- CP-element group 389: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1130_Sample/req
      -- 
    ack_2710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1127_inst_ack_1, ack => convTranspose_CP_39_elements(389)); -- 
    req_2718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(389), ack => WPIPE_Block1_start_1130_inst_req_0); -- 
    -- CP-element group 390:  transition  input  output  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	389 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	391 
    -- CP-element group 390:  members (6) 
      -- CP-element group 390: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1130_sample_completed_
      -- CP-element group 390: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1130_update_start_
      -- CP-element group 390: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1130_Sample/$exit
      -- CP-element group 390: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1130_Sample/ack
      -- CP-element group 390: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1130_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1130_Update/req
      -- 
    ack_2719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1130_inst_ack_0, ack => convTranspose_CP_39_elements(390)); -- 
    req_2723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(390), ack => WPIPE_Block1_start_1130_inst_req_1); -- 
    -- CP-element group 391:  transition  input  output  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	390 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	392 
    -- CP-element group 391:  members (6) 
      -- CP-element group 391: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1130_update_completed_
      -- CP-element group 391: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1130_Update/$exit
      -- CP-element group 391: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1130_Update/ack
      -- CP-element group 391: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1133_sample_start_
      -- CP-element group 391: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1133_Sample/$entry
      -- CP-element group 391: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1133_Sample/req
      -- 
    ack_2724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1130_inst_ack_1, ack => convTranspose_CP_39_elements(391)); -- 
    req_2732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(391), ack => WPIPE_Block1_start_1133_inst_req_0); -- 
    -- CP-element group 392:  transition  input  output  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	391 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	393 
    -- CP-element group 392:  members (6) 
      -- CP-element group 392: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1133_sample_completed_
      -- CP-element group 392: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1133_update_start_
      -- CP-element group 392: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1133_Sample/$exit
      -- CP-element group 392: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1133_Sample/ack
      -- CP-element group 392: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1133_Update/$entry
      -- CP-element group 392: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1133_Update/req
      -- 
    ack_2733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1133_inst_ack_0, ack => convTranspose_CP_39_elements(392)); -- 
    req_2737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(392), ack => WPIPE_Block1_start_1133_inst_req_1); -- 
    -- CP-element group 393:  transition  input  output  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	392 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	394 
    -- CP-element group 393:  members (6) 
      -- CP-element group 393: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1133_update_completed_
      -- CP-element group 393: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1133_Update/$exit
      -- CP-element group 393: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1133_Update/ack
      -- CP-element group 393: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1136_sample_start_
      -- CP-element group 393: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1136_Sample/$entry
      -- CP-element group 393: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1136_Sample/req
      -- 
    ack_2738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1133_inst_ack_1, ack => convTranspose_CP_39_elements(393)); -- 
    req_2746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(393), ack => WPIPE_Block1_start_1136_inst_req_0); -- 
    -- CP-element group 394:  transition  input  output  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	393 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	395 
    -- CP-element group 394:  members (6) 
      -- CP-element group 394: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1136_sample_completed_
      -- CP-element group 394: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1136_update_start_
      -- CP-element group 394: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1136_Sample/$exit
      -- CP-element group 394: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1136_Sample/ack
      -- CP-element group 394: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1136_Update/$entry
      -- CP-element group 394: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1136_Update/req
      -- 
    ack_2747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1136_inst_ack_0, ack => convTranspose_CP_39_elements(394)); -- 
    req_2751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(394), ack => WPIPE_Block1_start_1136_inst_req_1); -- 
    -- CP-element group 395:  transition  input  output  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	394 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	396 
    -- CP-element group 395:  members (6) 
      -- CP-element group 395: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1136_update_completed_
      -- CP-element group 395: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1136_Update/$exit
      -- CP-element group 395: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1136_Update/ack
      -- CP-element group 395: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1139_sample_start_
      -- CP-element group 395: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1139_Sample/$entry
      -- CP-element group 395: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1139_Sample/req
      -- 
    ack_2752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1136_inst_ack_1, ack => convTranspose_CP_39_elements(395)); -- 
    req_2760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(395), ack => WPIPE_Block1_start_1139_inst_req_0); -- 
    -- CP-element group 396:  transition  input  output  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	395 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	397 
    -- CP-element group 396:  members (6) 
      -- CP-element group 396: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1139_sample_completed_
      -- CP-element group 396: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1139_update_start_
      -- CP-element group 396: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1139_Sample/$exit
      -- CP-element group 396: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1139_Sample/ack
      -- CP-element group 396: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1139_Update/$entry
      -- CP-element group 396: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1139_Update/req
      -- 
    ack_2761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1139_inst_ack_0, ack => convTranspose_CP_39_elements(396)); -- 
    req_2765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(396), ack => WPIPE_Block1_start_1139_inst_req_1); -- 
    -- CP-element group 397:  transition  input  output  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	396 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	398 
    -- CP-element group 397:  members (6) 
      -- CP-element group 397: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1139_update_completed_
      -- CP-element group 397: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1139_Update/$exit
      -- CP-element group 397: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1139_Update/ack
      -- CP-element group 397: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1142_sample_start_
      -- CP-element group 397: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1142_Sample/$entry
      -- CP-element group 397: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1142_Sample/req
      -- 
    ack_2766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1139_inst_ack_1, ack => convTranspose_CP_39_elements(397)); -- 
    req_2774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(397), ack => WPIPE_Block1_start_1142_inst_req_0); -- 
    -- CP-element group 398:  transition  input  output  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	397 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	399 
    -- CP-element group 398:  members (6) 
      -- CP-element group 398: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1142_sample_completed_
      -- CP-element group 398: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1142_update_start_
      -- CP-element group 398: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1142_Sample/$exit
      -- CP-element group 398: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1142_Sample/ack
      -- CP-element group 398: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1142_Update/$entry
      -- CP-element group 398: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1142_Update/req
      -- 
    ack_2775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 398_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1142_inst_ack_0, ack => convTranspose_CP_39_elements(398)); -- 
    req_2779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(398), ack => WPIPE_Block1_start_1142_inst_req_1); -- 
    -- CP-element group 399:  transition  input  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	398 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	456 
    -- CP-element group 399:  members (3) 
      -- CP-element group 399: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1142_update_completed_
      -- CP-element group 399: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1142_Update/$exit
      -- CP-element group 399: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1142_Update/ack
      -- 
    ack_2780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1142_inst_ack_1, ack => convTranspose_CP_39_elements(399)); -- 
    -- CP-element group 400:  transition  input  output  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	535 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	401 
    -- CP-element group 400:  members (6) 
      -- CP-element group 400: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1145_sample_completed_
      -- CP-element group 400: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1145_update_start_
      -- CP-element group 400: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1145_Sample/$exit
      -- CP-element group 400: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1145_Sample/ack
      -- CP-element group 400: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1145_Update/$entry
      -- CP-element group 400: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1145_Update/req
      -- 
    ack_2789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1145_inst_ack_0, ack => convTranspose_CP_39_elements(400)); -- 
    req_2793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(400), ack => WPIPE_Block2_start_1145_inst_req_1); -- 
    -- CP-element group 401:  transition  input  output  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	400 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	402 
    -- CP-element group 401:  members (6) 
      -- CP-element group 401: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1145_update_completed_
      -- CP-element group 401: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1145_Update/$exit
      -- CP-element group 401: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1145_Update/ack
      -- CP-element group 401: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1148_sample_start_
      -- CP-element group 401: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1148_Sample/$entry
      -- CP-element group 401: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1148_Sample/req
      -- 
    ack_2794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1145_inst_ack_1, ack => convTranspose_CP_39_elements(401)); -- 
    req_2802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(401), ack => WPIPE_Block2_start_1148_inst_req_0); -- 
    -- CP-element group 402:  transition  input  output  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	401 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	403 
    -- CP-element group 402:  members (6) 
      -- CP-element group 402: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1148_sample_completed_
      -- CP-element group 402: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1148_update_start_
      -- CP-element group 402: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1148_Sample/$exit
      -- CP-element group 402: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1148_Sample/ack
      -- CP-element group 402: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1148_Update/$entry
      -- CP-element group 402: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1148_Update/req
      -- 
    ack_2803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 402_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1148_inst_ack_0, ack => convTranspose_CP_39_elements(402)); -- 
    req_2807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(402), ack => WPIPE_Block2_start_1148_inst_req_1); -- 
    -- CP-element group 403:  transition  input  output  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	402 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	404 
    -- CP-element group 403:  members (6) 
      -- CP-element group 403: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1148_update_completed_
      -- CP-element group 403: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1148_Update/$exit
      -- CP-element group 403: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1148_Update/ack
      -- CP-element group 403: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1151_sample_start_
      -- CP-element group 403: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1151_Sample/$entry
      -- CP-element group 403: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1151_Sample/req
      -- 
    ack_2808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1148_inst_ack_1, ack => convTranspose_CP_39_elements(403)); -- 
    req_2816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(403), ack => WPIPE_Block2_start_1151_inst_req_0); -- 
    -- CP-element group 404:  transition  input  output  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	403 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	405 
    -- CP-element group 404:  members (6) 
      -- CP-element group 404: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1151_sample_completed_
      -- CP-element group 404: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1151_update_start_
      -- CP-element group 404: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1151_Sample/$exit
      -- CP-element group 404: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1151_Sample/ack
      -- CP-element group 404: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1151_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1151_Update/req
      -- 
    ack_2817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1151_inst_ack_0, ack => convTranspose_CP_39_elements(404)); -- 
    req_2821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => WPIPE_Block2_start_1151_inst_req_1); -- 
    -- CP-element group 405:  transition  input  output  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	404 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	406 
    -- CP-element group 405:  members (6) 
      -- CP-element group 405: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1151_update_completed_
      -- CP-element group 405: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1151_Update/$exit
      -- CP-element group 405: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1151_Update/ack
      -- CP-element group 405: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1154_sample_start_
      -- CP-element group 405: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1154_Sample/$entry
      -- CP-element group 405: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1154_Sample/req
      -- 
    ack_2822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 405_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1151_inst_ack_1, ack => convTranspose_CP_39_elements(405)); -- 
    req_2830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(405), ack => WPIPE_Block2_start_1154_inst_req_0); -- 
    -- CP-element group 406:  transition  input  output  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	405 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	407 
    -- CP-element group 406:  members (6) 
      -- CP-element group 406: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1154_sample_completed_
      -- CP-element group 406: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1154_update_start_
      -- CP-element group 406: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1154_Sample/$exit
      -- CP-element group 406: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1154_Sample/ack
      -- CP-element group 406: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1154_Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1154_Update/req
      -- 
    ack_2831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 406_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1154_inst_ack_0, ack => convTranspose_CP_39_elements(406)); -- 
    req_2835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(406), ack => WPIPE_Block2_start_1154_inst_req_1); -- 
    -- CP-element group 407:  transition  input  output  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	406 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	408 
    -- CP-element group 407:  members (6) 
      -- CP-element group 407: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1154_update_completed_
      -- CP-element group 407: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1154_Update/$exit
      -- CP-element group 407: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1154_Update/ack
      -- CP-element group 407: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1157_sample_start_
      -- CP-element group 407: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1157_Sample/$entry
      -- CP-element group 407: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1157_Sample/req
      -- 
    ack_2836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1154_inst_ack_1, ack => convTranspose_CP_39_elements(407)); -- 
    req_2844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(407), ack => WPIPE_Block2_start_1157_inst_req_0); -- 
    -- CP-element group 408:  transition  input  output  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	407 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	409 
    -- CP-element group 408:  members (6) 
      -- CP-element group 408: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1157_sample_completed_
      -- CP-element group 408: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1157_update_start_
      -- CP-element group 408: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1157_Sample/$exit
      -- CP-element group 408: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1157_Sample/ack
      -- CP-element group 408: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1157_Update/$entry
      -- CP-element group 408: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1157_Update/req
      -- 
    ack_2845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 408_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1157_inst_ack_0, ack => convTranspose_CP_39_elements(408)); -- 
    req_2849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(408), ack => WPIPE_Block2_start_1157_inst_req_1); -- 
    -- CP-element group 409:  transition  input  output  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	408 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	410 
    -- CP-element group 409:  members (6) 
      -- CP-element group 409: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1157_update_completed_
      -- CP-element group 409: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1157_Update/$exit
      -- CP-element group 409: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1157_Update/ack
      -- CP-element group 409: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1160_sample_start_
      -- CP-element group 409: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1160_Sample/$entry
      -- CP-element group 409: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1160_Sample/req
      -- 
    ack_2850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 409_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1157_inst_ack_1, ack => convTranspose_CP_39_elements(409)); -- 
    req_2858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(409), ack => WPIPE_Block2_start_1160_inst_req_0); -- 
    -- CP-element group 410:  transition  input  output  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	409 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	411 
    -- CP-element group 410:  members (6) 
      -- CP-element group 410: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1160_sample_completed_
      -- CP-element group 410: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1160_update_start_
      -- CP-element group 410: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1160_Sample/$exit
      -- CP-element group 410: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1160_Sample/ack
      -- CP-element group 410: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1160_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1160_Update/req
      -- 
    ack_2859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1160_inst_ack_0, ack => convTranspose_CP_39_elements(410)); -- 
    req_2863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => WPIPE_Block2_start_1160_inst_req_1); -- 
    -- CP-element group 411:  transition  input  output  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	410 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	412 
    -- CP-element group 411:  members (6) 
      -- CP-element group 411: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1160_update_completed_
      -- CP-element group 411: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1160_Update/$exit
      -- CP-element group 411: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1160_Update/ack
      -- CP-element group 411: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1163_sample_start_
      -- CP-element group 411: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1163_Sample/$entry
      -- CP-element group 411: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1163_Sample/req
      -- 
    ack_2864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 411_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1160_inst_ack_1, ack => convTranspose_CP_39_elements(411)); -- 
    req_2872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(411), ack => WPIPE_Block2_start_1163_inst_req_0); -- 
    -- CP-element group 412:  transition  input  output  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	411 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	413 
    -- CP-element group 412:  members (6) 
      -- CP-element group 412: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1163_sample_completed_
      -- CP-element group 412: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1163_update_start_
      -- CP-element group 412: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1163_Sample/$exit
      -- CP-element group 412: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1163_Sample/ack
      -- CP-element group 412: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1163_Update/$entry
      -- CP-element group 412: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1163_Update/req
      -- 
    ack_2873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1163_inst_ack_0, ack => convTranspose_CP_39_elements(412)); -- 
    req_2877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(412), ack => WPIPE_Block2_start_1163_inst_req_1); -- 
    -- CP-element group 413:  transition  input  output  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	412 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	414 
    -- CP-element group 413:  members (6) 
      -- CP-element group 413: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1163_update_completed_
      -- CP-element group 413: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1163_Update/$exit
      -- CP-element group 413: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1163_Update/ack
      -- CP-element group 413: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1166_sample_start_
      -- CP-element group 413: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1166_Sample/$entry
      -- CP-element group 413: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1166_Sample/req
      -- 
    ack_2878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1163_inst_ack_1, ack => convTranspose_CP_39_elements(413)); -- 
    req_2886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(413), ack => WPIPE_Block2_start_1166_inst_req_0); -- 
    -- CP-element group 414:  transition  input  output  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	413 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	415 
    -- CP-element group 414:  members (6) 
      -- CP-element group 414: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1166_sample_completed_
      -- CP-element group 414: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1166_update_start_
      -- CP-element group 414: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1166_Sample/$exit
      -- CP-element group 414: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1166_Sample/ack
      -- CP-element group 414: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1166_Update/$entry
      -- CP-element group 414: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1166_Update/req
      -- 
    ack_2887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 414_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1166_inst_ack_0, ack => convTranspose_CP_39_elements(414)); -- 
    req_2891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(414), ack => WPIPE_Block2_start_1166_inst_req_1); -- 
    -- CP-element group 415:  transition  input  output  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	414 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	416 
    -- CP-element group 415:  members (6) 
      -- CP-element group 415: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1166_update_completed_
      -- CP-element group 415: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1166_Update/$exit
      -- CP-element group 415: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1166_Update/ack
      -- CP-element group 415: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1169_sample_start_
      -- CP-element group 415: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1169_Sample/$entry
      -- CP-element group 415: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1169_Sample/req
      -- 
    ack_2892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 415_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1166_inst_ack_1, ack => convTranspose_CP_39_elements(415)); -- 
    req_2900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(415), ack => WPIPE_Block2_start_1169_inst_req_0); -- 
    -- CP-element group 416:  transition  input  output  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	415 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	417 
    -- CP-element group 416:  members (6) 
      -- CP-element group 416: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1169_sample_completed_
      -- CP-element group 416: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1169_update_start_
      -- CP-element group 416: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1169_Sample/$exit
      -- CP-element group 416: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1169_Sample/ack
      -- CP-element group 416: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1169_Update/$entry
      -- CP-element group 416: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1169_Update/req
      -- 
    ack_2901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1169_inst_ack_0, ack => convTranspose_CP_39_elements(416)); -- 
    req_2905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(416), ack => WPIPE_Block2_start_1169_inst_req_1); -- 
    -- CP-element group 417:  transition  input  output  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	416 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	418 
    -- CP-element group 417:  members (6) 
      -- CP-element group 417: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1169_update_completed_
      -- CP-element group 417: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1169_Update/$exit
      -- CP-element group 417: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1169_Update/ack
      -- CP-element group 417: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1172_sample_start_
      -- CP-element group 417: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1172_Sample/$entry
      -- CP-element group 417: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1172_Sample/req
      -- 
    ack_2906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1169_inst_ack_1, ack => convTranspose_CP_39_elements(417)); -- 
    req_2914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(417), ack => WPIPE_Block2_start_1172_inst_req_0); -- 
    -- CP-element group 418:  transition  input  output  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	417 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	419 
    -- CP-element group 418:  members (6) 
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1172_sample_completed_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1172_update_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1172_Sample/$exit
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1172_Sample/ack
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1172_Update/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1172_Update/req
      -- 
    ack_2915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 418_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1172_inst_ack_0, ack => convTranspose_CP_39_elements(418)); -- 
    req_2919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => WPIPE_Block2_start_1172_inst_req_1); -- 
    -- CP-element group 419:  transition  input  output  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	418 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	420 
    -- CP-element group 419:  members (6) 
      -- CP-element group 419: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1172_update_completed_
      -- CP-element group 419: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1172_Update/$exit
      -- CP-element group 419: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1172_Update/ack
      -- CP-element group 419: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1175_sample_start_
      -- CP-element group 419: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1175_Sample/$entry
      -- CP-element group 419: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1175_Sample/req
      -- 
    ack_2920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1172_inst_ack_1, ack => convTranspose_CP_39_elements(419)); -- 
    req_2928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(419), ack => WPIPE_Block2_start_1175_inst_req_0); -- 
    -- CP-element group 420:  transition  input  output  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	419 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	421 
    -- CP-element group 420:  members (6) 
      -- CP-element group 420: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1175_sample_completed_
      -- CP-element group 420: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1175_update_start_
      -- CP-element group 420: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1175_Sample/$exit
      -- CP-element group 420: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1175_Sample/ack
      -- CP-element group 420: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1175_Update/$entry
      -- CP-element group 420: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1175_Update/req
      -- 
    ack_2929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1175_inst_ack_0, ack => convTranspose_CP_39_elements(420)); -- 
    req_2933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(420), ack => WPIPE_Block2_start_1175_inst_req_1); -- 
    -- CP-element group 421:  transition  input  output  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	420 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	422 
    -- CP-element group 421:  members (6) 
      -- CP-element group 421: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1175_update_completed_
      -- CP-element group 421: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1175_Update/$exit
      -- CP-element group 421: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1175_Update/ack
      -- CP-element group 421: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1178_sample_start_
      -- CP-element group 421: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1178_Sample/$entry
      -- CP-element group 421: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1178_Sample/req
      -- 
    ack_2934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1175_inst_ack_1, ack => convTranspose_CP_39_elements(421)); -- 
    req_2942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(421), ack => WPIPE_Block2_start_1178_inst_req_0); -- 
    -- CP-element group 422:  transition  input  output  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	421 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	423 
    -- CP-element group 422:  members (6) 
      -- CP-element group 422: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1178_sample_completed_
      -- CP-element group 422: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1178_update_start_
      -- CP-element group 422: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1178_Sample/$exit
      -- CP-element group 422: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1178_Sample/ack
      -- CP-element group 422: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1178_Update/$entry
      -- CP-element group 422: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1178_Update/req
      -- 
    ack_2943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 422_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1178_inst_ack_0, ack => convTranspose_CP_39_elements(422)); -- 
    req_2947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(422), ack => WPIPE_Block2_start_1178_inst_req_1); -- 
    -- CP-element group 423:  transition  input  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	422 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	456 
    -- CP-element group 423:  members (3) 
      -- CP-element group 423: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1178_update_completed_
      -- CP-element group 423: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1178_Update/$exit
      -- CP-element group 423: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1178_Update/ack
      -- 
    ack_2948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 423_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1178_inst_ack_1, ack => convTranspose_CP_39_elements(423)); -- 
    -- CP-element group 424:  transition  input  output  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	535 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	425 
    -- CP-element group 424:  members (6) 
      -- CP-element group 424: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1181_sample_completed_
      -- CP-element group 424: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1181_update_start_
      -- CP-element group 424: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1181_Sample/$exit
      -- CP-element group 424: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1181_Sample/ack
      -- CP-element group 424: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1181_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1181_Update/req
      -- 
    ack_2957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1181_inst_ack_0, ack => convTranspose_CP_39_elements(424)); -- 
    req_2961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => WPIPE_Block3_start_1181_inst_req_1); -- 
    -- CP-element group 425:  transition  input  output  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	424 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	426 
    -- CP-element group 425:  members (6) 
      -- CP-element group 425: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1181_update_completed_
      -- CP-element group 425: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1181_Update/$exit
      -- CP-element group 425: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1181_Update/ack
      -- CP-element group 425: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1184_sample_start_
      -- CP-element group 425: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1184_Sample/$entry
      -- CP-element group 425: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1184_Sample/req
      -- 
    ack_2962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1181_inst_ack_1, ack => convTranspose_CP_39_elements(425)); -- 
    req_2970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(425), ack => WPIPE_Block3_start_1184_inst_req_0); -- 
    -- CP-element group 426:  transition  input  output  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	425 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	427 
    -- CP-element group 426:  members (6) 
      -- CP-element group 426: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1184_sample_completed_
      -- CP-element group 426: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1184_update_start_
      -- CP-element group 426: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1184_Sample/$exit
      -- CP-element group 426: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1184_Sample/ack
      -- CP-element group 426: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1184_Update/$entry
      -- CP-element group 426: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1184_Update/req
      -- 
    ack_2971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 426_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1184_inst_ack_0, ack => convTranspose_CP_39_elements(426)); -- 
    req_2975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(426), ack => WPIPE_Block3_start_1184_inst_req_1); -- 
    -- CP-element group 427:  transition  input  output  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	426 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	428 
    -- CP-element group 427:  members (6) 
      -- CP-element group 427: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1184_update_completed_
      -- CP-element group 427: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1184_Update/$exit
      -- CP-element group 427: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1184_Update/ack
      -- CP-element group 427: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1187_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1187_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1187_Sample/req
      -- 
    ack_2976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 427_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1184_inst_ack_1, ack => convTranspose_CP_39_elements(427)); -- 
    req_2984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(427), ack => WPIPE_Block3_start_1187_inst_req_0); -- 
    -- CP-element group 428:  transition  input  output  bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	427 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	429 
    -- CP-element group 428:  members (6) 
      -- CP-element group 428: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1187_sample_completed_
      -- CP-element group 428: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1187_update_start_
      -- CP-element group 428: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1187_Sample/$exit
      -- CP-element group 428: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1187_Sample/ack
      -- CP-element group 428: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1187_Update/$entry
      -- CP-element group 428: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1187_Update/req
      -- 
    ack_2985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1187_inst_ack_0, ack => convTranspose_CP_39_elements(428)); -- 
    req_2989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(428), ack => WPIPE_Block3_start_1187_inst_req_1); -- 
    -- CP-element group 429:  transition  input  output  bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	428 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	430 
    -- CP-element group 429:  members (6) 
      -- CP-element group 429: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1187_update_completed_
      -- CP-element group 429: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1187_Update/$exit
      -- CP-element group 429: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1187_Update/ack
      -- CP-element group 429: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1190_sample_start_
      -- CP-element group 429: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1190_Sample/$entry
      -- CP-element group 429: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1190_Sample/req
      -- 
    ack_2990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1187_inst_ack_1, ack => convTranspose_CP_39_elements(429)); -- 
    req_2998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(429), ack => WPIPE_Block3_start_1190_inst_req_0); -- 
    -- CP-element group 430:  transition  input  output  bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	429 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	431 
    -- CP-element group 430:  members (6) 
      -- CP-element group 430: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1190_sample_completed_
      -- CP-element group 430: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1190_update_start_
      -- CP-element group 430: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1190_Sample/$exit
      -- CP-element group 430: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1190_Sample/ack
      -- CP-element group 430: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1190_Update/$entry
      -- CP-element group 430: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1190_Update/req
      -- 
    ack_2999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 430_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1190_inst_ack_0, ack => convTranspose_CP_39_elements(430)); -- 
    req_3003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(430), ack => WPIPE_Block3_start_1190_inst_req_1); -- 
    -- CP-element group 431:  transition  input  output  bypass 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	430 
    -- CP-element group 431: successors 
    -- CP-element group 431: 	432 
    -- CP-element group 431:  members (6) 
      -- CP-element group 431: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1190_update_completed_
      -- CP-element group 431: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1190_Update/$exit
      -- CP-element group 431: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1190_Update/ack
      -- CP-element group 431: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1193_sample_start_
      -- CP-element group 431: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1193_Sample/$entry
      -- CP-element group 431: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1193_Sample/req
      -- 
    ack_3004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 431_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1190_inst_ack_1, ack => convTranspose_CP_39_elements(431)); -- 
    req_3012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(431), ack => WPIPE_Block3_start_1193_inst_req_0); -- 
    -- CP-element group 432:  transition  input  output  bypass 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	431 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	433 
    -- CP-element group 432:  members (6) 
      -- CP-element group 432: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1193_Update/req
      -- CP-element group 432: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1193_Update/$entry
      -- CP-element group 432: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1193_sample_completed_
      -- CP-element group 432: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1193_update_start_
      -- CP-element group 432: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1193_Sample/$exit
      -- CP-element group 432: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1193_Sample/ack
      -- 
    ack_3013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1193_inst_ack_0, ack => convTranspose_CP_39_elements(432)); -- 
    req_3017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(432), ack => WPIPE_Block3_start_1193_inst_req_1); -- 
    -- CP-element group 433:  transition  input  output  bypass 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	432 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	434 
    -- CP-element group 433:  members (6) 
      -- CP-element group 433: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1196_Sample/$entry
      -- CP-element group 433: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1196_Sample/req
      -- CP-element group 433: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1196_sample_start_
      -- CP-element group 433: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1193_Update/ack
      -- CP-element group 433: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1193_Update/$exit
      -- CP-element group 433: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1193_update_completed_
      -- 
    ack_3018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1193_inst_ack_1, ack => convTranspose_CP_39_elements(433)); -- 
    req_3026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(433), ack => WPIPE_Block3_start_1196_inst_req_0); -- 
    -- CP-element group 434:  transition  input  output  bypass 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	433 
    -- CP-element group 434: successors 
    -- CP-element group 434: 	435 
    -- CP-element group 434:  members (6) 
      -- CP-element group 434: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1196_Update/req
      -- CP-element group 434: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1196_update_start_
      -- CP-element group 434: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1196_Sample/$exit
      -- CP-element group 434: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1196_sample_completed_
      -- CP-element group 434: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1196_Update/$entry
      -- CP-element group 434: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1196_Sample/ack
      -- 
    ack_3027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 434_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1196_inst_ack_0, ack => convTranspose_CP_39_elements(434)); -- 
    req_3031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(434), ack => WPIPE_Block3_start_1196_inst_req_1); -- 
    -- CP-element group 435:  transition  input  output  bypass 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	434 
    -- CP-element group 435: successors 
    -- CP-element group 435: 	436 
    -- CP-element group 435:  members (6) 
      -- CP-element group 435: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1196_Update/ack
      -- CP-element group 435: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1199_sample_start_
      -- CP-element group 435: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1196_update_completed_
      -- CP-element group 435: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1199_Sample/$entry
      -- CP-element group 435: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1196_Update/$exit
      -- CP-element group 435: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1199_Sample/req
      -- 
    ack_3032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1196_inst_ack_1, ack => convTranspose_CP_39_elements(435)); -- 
    req_3040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(435), ack => WPIPE_Block3_start_1199_inst_req_0); -- 
    -- CP-element group 436:  transition  input  output  bypass 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	435 
    -- CP-element group 436: successors 
    -- CP-element group 436: 	437 
    -- CP-element group 436:  members (6) 
      -- CP-element group 436: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1199_sample_completed_
      -- CP-element group 436: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1199_update_start_
      -- CP-element group 436: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1199_Sample/$exit
      -- CP-element group 436: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1199_Update/req
      -- CP-element group 436: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1199_Update/$entry
      -- CP-element group 436: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1199_Sample/ack
      -- 
    ack_3041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1199_inst_ack_0, ack => convTranspose_CP_39_elements(436)); -- 
    req_3045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(436), ack => WPIPE_Block3_start_1199_inst_req_1); -- 
    -- CP-element group 437:  transition  input  output  bypass 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	436 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	438 
    -- CP-element group 437:  members (6) 
      -- CP-element group 437: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1199_update_completed_
      -- CP-element group 437: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1202_Sample/req
      -- CP-element group 437: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1202_Sample/$entry
      -- CP-element group 437: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1202_sample_start_
      -- CP-element group 437: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1199_Update/ack
      -- CP-element group 437: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1199_Update/$exit
      -- 
    ack_3046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 437_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1199_inst_ack_1, ack => convTranspose_CP_39_elements(437)); -- 
    req_3054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(437), ack => WPIPE_Block3_start_1202_inst_req_0); -- 
    -- CP-element group 438:  transition  input  output  bypass 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	437 
    -- CP-element group 438: successors 
    -- CP-element group 438: 	439 
    -- CP-element group 438:  members (6) 
      -- CP-element group 438: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1202_Update/req
      -- CP-element group 438: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1202_Update/$entry
      -- CP-element group 438: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1202_Sample/ack
      -- CP-element group 438: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1202_Sample/$exit
      -- CP-element group 438: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1202_update_start_
      -- CP-element group 438: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1202_sample_completed_
      -- 
    ack_3055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 438_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1202_inst_ack_0, ack => convTranspose_CP_39_elements(438)); -- 
    req_3059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(438), ack => WPIPE_Block3_start_1202_inst_req_1); -- 
    -- CP-element group 439:  transition  input  output  bypass 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	438 
    -- CP-element group 439: successors 
    -- CP-element group 439: 	440 
    -- CP-element group 439:  members (6) 
      -- CP-element group 439: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1205_Sample/req
      -- CP-element group 439: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1205_Sample/$entry
      -- CP-element group 439: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1205_sample_start_
      -- CP-element group 439: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1202_Update/ack
      -- CP-element group 439: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1202_Update/$exit
      -- CP-element group 439: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1202_update_completed_
      -- 
    ack_3060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 439_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1202_inst_ack_1, ack => convTranspose_CP_39_elements(439)); -- 
    req_3068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(439), ack => WPIPE_Block3_start_1205_inst_req_0); -- 
    -- CP-element group 440:  transition  input  output  bypass 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	439 
    -- CP-element group 440: successors 
    -- CP-element group 440: 	441 
    -- CP-element group 440:  members (6) 
      -- CP-element group 440: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1205_Update/req
      -- CP-element group 440: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1205_Update/$entry
      -- CP-element group 440: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1205_Sample/ack
      -- CP-element group 440: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1205_Sample/$exit
      -- CP-element group 440: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1205_update_start_
      -- CP-element group 440: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1205_sample_completed_
      -- 
    ack_3069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 440_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1205_inst_ack_0, ack => convTranspose_CP_39_elements(440)); -- 
    req_3073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(440), ack => WPIPE_Block3_start_1205_inst_req_1); -- 
    -- CP-element group 441:  transition  input  output  bypass 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	440 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	442 
    -- CP-element group 441:  members (6) 
      -- CP-element group 441: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1208_Sample/req
      -- CP-element group 441: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1208_Sample/$entry
      -- CP-element group 441: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1208_sample_start_
      -- CP-element group 441: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1205_Update/ack
      -- CP-element group 441: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1205_Update/$exit
      -- CP-element group 441: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1205_update_completed_
      -- 
    ack_3074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 441_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1205_inst_ack_1, ack => convTranspose_CP_39_elements(441)); -- 
    req_3082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(441), ack => WPIPE_Block3_start_1208_inst_req_0); -- 
    -- CP-element group 442:  transition  input  output  bypass 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	441 
    -- CP-element group 442: successors 
    -- CP-element group 442: 	443 
    -- CP-element group 442:  members (6) 
      -- CP-element group 442: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1208_update_start_
      -- CP-element group 442: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1208_sample_completed_
      -- CP-element group 442: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1208_Update/$entry
      -- CP-element group 442: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1208_Sample/$exit
      -- CP-element group 442: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1208_Sample/ack
      -- CP-element group 442: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1208_Update/req
      -- 
    ack_3083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 442_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1208_inst_ack_0, ack => convTranspose_CP_39_elements(442)); -- 
    req_3087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(442), ack => WPIPE_Block3_start_1208_inst_req_1); -- 
    -- CP-element group 443:  transition  input  output  bypass 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	442 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	444 
    -- CP-element group 443:  members (6) 
      -- CP-element group 443: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1208_update_completed_
      -- CP-element group 443: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1208_Update/$exit
      -- CP-element group 443: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1208_Update/ack
      -- CP-element group 443: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1211_sample_start_
      -- CP-element group 443: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1211_Sample/$entry
      -- CP-element group 443: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1211_Sample/req
      -- 
    ack_3088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 443_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1208_inst_ack_1, ack => convTranspose_CP_39_elements(443)); -- 
    req_3096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(443), ack => WPIPE_Block3_start_1211_inst_req_0); -- 
    -- CP-element group 444:  transition  input  output  bypass 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	443 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	445 
    -- CP-element group 444:  members (6) 
      -- CP-element group 444: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1211_Update/req
      -- CP-element group 444: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1211_sample_completed_
      -- CP-element group 444: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1211_update_start_
      -- CP-element group 444: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1211_Sample/$exit
      -- CP-element group 444: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1211_Update/$entry
      -- CP-element group 444: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1211_Sample/ack
      -- 
    ack_3097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1211_inst_ack_0, ack => convTranspose_CP_39_elements(444)); -- 
    req_3101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(444), ack => WPIPE_Block3_start_1211_inst_req_1); -- 
    -- CP-element group 445:  transition  input  output  bypass 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	444 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	446 
    -- CP-element group 445:  members (6) 
      -- CP-element group 445: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1211_Update/ack
      -- CP-element group 445: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1214_sample_start_
      -- CP-element group 445: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1211_update_completed_
      -- CP-element group 445: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1211_Update/$exit
      -- CP-element group 445: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1214_Sample/req
      -- CP-element group 445: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1214_Sample/$entry
      -- 
    ack_3102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 445_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1211_inst_ack_1, ack => convTranspose_CP_39_elements(445)); -- 
    req_3110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(445), ack => WPIPE_Block3_start_1214_inst_req_0); -- 
    -- CP-element group 446:  transition  input  output  bypass 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	445 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	447 
    -- CP-element group 446:  members (6) 
      -- CP-element group 446: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1214_sample_completed_
      -- CP-element group 446: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1214_update_start_
      -- CP-element group 446: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1214_Update/req
      -- CP-element group 446: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1214_Update/$entry
      -- CP-element group 446: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1214_Sample/ack
      -- CP-element group 446: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1214_Sample/$exit
      -- 
    ack_3111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 446_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1214_inst_ack_0, ack => convTranspose_CP_39_elements(446)); -- 
    req_3115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(446), ack => WPIPE_Block3_start_1214_inst_req_1); -- 
    -- CP-element group 447:  transition  input  bypass 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	446 
    -- CP-element group 447: successors 
    -- CP-element group 447: 	456 
    -- CP-element group 447:  members (3) 
      -- CP-element group 447: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1214_update_completed_
      -- CP-element group 447: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1214_Update/ack
      -- CP-element group 447: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1214_Update/$exit
      -- 
    ack_3116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1214_inst_ack_1, ack => convTranspose_CP_39_elements(447)); -- 
    -- CP-element group 448:  transition  input  output  bypass 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	535 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	449 
    -- CP-element group 448:  members (6) 
      -- CP-element group 448: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block0_done_1218_Update/cr
      -- CP-element group 448: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block0_done_1218_Update/$entry
      -- CP-element group 448: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block0_done_1218_Sample/ra
      -- CP-element group 448: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block0_done_1218_Sample/$exit
      -- CP-element group 448: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block0_done_1218_update_start_
      -- CP-element group 448: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block0_done_1218_sample_completed_
      -- 
    ra_3125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 448_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1218_inst_ack_0, ack => convTranspose_CP_39_elements(448)); -- 
    cr_3129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(448), ack => RPIPE_Block0_done_1218_inst_req_1); -- 
    -- CP-element group 449:  transition  input  bypass 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	448 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	456 
    -- CP-element group 449:  members (3) 
      -- CP-element group 449: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block0_done_1218_Update/ca
      -- CP-element group 449: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block0_done_1218_Update/$exit
      -- CP-element group 449: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block0_done_1218_update_completed_
      -- 
    ca_3130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 449_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1218_inst_ack_1, ack => convTranspose_CP_39_elements(449)); -- 
    -- CP-element group 450:  transition  input  output  bypass 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	535 
    -- CP-element group 450: successors 
    -- CP-element group 450: 	451 
    -- CP-element group 450:  members (6) 
      -- CP-element group 450: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block1_done_1221_Update/cr
      -- CP-element group 450: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block1_done_1221_Update/$entry
      -- CP-element group 450: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block1_done_1221_Sample/ra
      -- CP-element group 450: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block1_done_1221_Sample/$exit
      -- CP-element group 450: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block1_done_1221_update_start_
      -- CP-element group 450: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block1_done_1221_sample_completed_
      -- 
    ra_3139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 450_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1221_inst_ack_0, ack => convTranspose_CP_39_elements(450)); -- 
    cr_3143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(450), ack => RPIPE_Block1_done_1221_inst_req_1); -- 
    -- CP-element group 451:  transition  input  bypass 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	450 
    -- CP-element group 451: successors 
    -- CP-element group 451: 	456 
    -- CP-element group 451:  members (3) 
      -- CP-element group 451: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block1_done_1221_Update/ca
      -- CP-element group 451: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block1_done_1221_Update/$exit
      -- CP-element group 451: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block1_done_1221_update_completed_
      -- 
    ca_3144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 451_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1221_inst_ack_1, ack => convTranspose_CP_39_elements(451)); -- 
    -- CP-element group 452:  transition  input  output  bypass 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	535 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	453 
    -- CP-element group 452:  members (6) 
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block2_done_1224_Update/cr
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block2_done_1224_Update/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block2_done_1224_Sample/ra
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block2_done_1224_Sample/$exit
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block2_done_1224_update_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block2_done_1224_sample_completed_
      -- 
    ra_3153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 452_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1224_inst_ack_0, ack => convTranspose_CP_39_elements(452)); -- 
    cr_3157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => RPIPE_Block2_done_1224_inst_req_1); -- 
    -- CP-element group 453:  transition  input  bypass 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	452 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	456 
    -- CP-element group 453:  members (3) 
      -- CP-element group 453: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block2_done_1224_Update/ca
      -- CP-element group 453: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block2_done_1224_Update/$exit
      -- CP-element group 453: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block2_done_1224_update_completed_
      -- 
    ca_3158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 453_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1224_inst_ack_1, ack => convTranspose_CP_39_elements(453)); -- 
    -- CP-element group 454:  transition  input  output  bypass 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	535 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	455 
    -- CP-element group 454:  members (6) 
      -- CP-element group 454: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block3_done_1227_Update/$entry
      -- CP-element group 454: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block3_done_1227_Sample/ra
      -- CP-element group 454: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block3_done_1227_Sample/$exit
      -- CP-element group 454: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block3_done_1227_Update/cr
      -- CP-element group 454: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block3_done_1227_update_start_
      -- CP-element group 454: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block3_done_1227_sample_completed_
      -- 
    ra_3167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 454_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1227_inst_ack_0, ack => convTranspose_CP_39_elements(454)); -- 
    cr_3171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(454), ack => RPIPE_Block3_done_1227_inst_req_1); -- 
    -- CP-element group 455:  transition  input  bypass 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	454 
    -- CP-element group 455: successors 
    -- CP-element group 455: 	456 
    -- CP-element group 455:  members (3) 
      -- CP-element group 455: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block3_done_1227_update_completed_
      -- CP-element group 455: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block3_done_1227_Update/$exit
      -- CP-element group 455: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block3_done_1227_Update/ca
      -- 
    ca_3172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 455_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1227_inst_ack_1, ack => convTranspose_CP_39_elements(455)); -- 
    -- CP-element group 456:  join  fork  transition  place  output  bypass 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	351 
    -- CP-element group 456: 	375 
    -- CP-element group 456: 	423 
    -- CP-element group 456: 	447 
    -- CP-element group 456: 	449 
    -- CP-element group 456: 	451 
    -- CP-element group 456: 	453 
    -- CP-element group 456: 	455 
    -- CP-element group 456: 	399 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	457 
    -- CP-element group 456: 	458 
    -- CP-element group 456: 	460 
    -- CP-element group 456:  members (13) 
      -- CP-element group 456: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228__exit__
      -- CP-element group 456: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244__entry__
      -- CP-element group 456: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/type_cast_1235_update_start_
      -- CP-element group 456: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/type_cast_1235_Update/$entry
      -- CP-element group 456: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/call_stmt_1231_Sample/$entry
      -- CP-element group 456: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/call_stmt_1231_sample_start_
      -- CP-element group 456: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/call_stmt_1231_update_start_
      -- CP-element group 456: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/type_cast_1235_Update/cr
      -- CP-element group 456: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/call_stmt_1231_Sample/crr
      -- CP-element group 456: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/call_stmt_1231_Update/$entry
      -- CP-element group 456: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/call_stmt_1231_Update/ccr
      -- CP-element group 456: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/$exit
      -- CP-element group 456: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/$entry
      -- 
    cr_3202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(456), ack => type_cast_1235_inst_req_1); -- 
    crr_3183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(456), ack => call_stmt_1231_call_req_0); -- 
    ccr_3188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(456), ack => call_stmt_1231_call_req_1); -- 
    convTranspose_cp_element_group_456: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_456"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(351) & convTranspose_CP_39_elements(375) & convTranspose_CP_39_elements(423) & convTranspose_CP_39_elements(447) & convTranspose_CP_39_elements(449) & convTranspose_CP_39_elements(451) & convTranspose_CP_39_elements(453) & convTranspose_CP_39_elements(455) & convTranspose_CP_39_elements(399);
      gj_convTranspose_cp_element_group_456 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(456), clk => clk, reset => reset); --
    end block;
    -- CP-element group 457:  transition  input  bypass 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	456 
    -- CP-element group 457: successors 
    -- CP-element group 457:  members (3) 
      -- CP-element group 457: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/call_stmt_1231_Sample/$exit
      -- CP-element group 457: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/call_stmt_1231_sample_completed_
      -- CP-element group 457: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/call_stmt_1231_Sample/cra
      -- 
    cra_3184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 457_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1231_call_ack_0, ack => convTranspose_CP_39_elements(457)); -- 
    -- CP-element group 458:  transition  input  output  bypass 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	456 
    -- CP-element group 458: successors 
    -- CP-element group 458: 	459 
    -- CP-element group 458:  members (6) 
      -- CP-element group 458: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/type_cast_1235_Sample/rr
      -- CP-element group 458: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/call_stmt_1231_update_completed_
      -- CP-element group 458: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/call_stmt_1231_Update/$exit
      -- CP-element group 458: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/call_stmt_1231_Update/cca
      -- CP-element group 458: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/type_cast_1235_sample_start_
      -- CP-element group 458: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/type_cast_1235_Sample/$entry
      -- 
    cca_3189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 458_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1231_call_ack_1, ack => convTranspose_CP_39_elements(458)); -- 
    rr_3197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(458), ack => type_cast_1235_inst_req_0); -- 
    -- CP-element group 459:  transition  input  bypass 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	458 
    -- CP-element group 459: successors 
    -- CP-element group 459:  members (3) 
      -- CP-element group 459: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/type_cast_1235_Sample/ra
      -- CP-element group 459: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/type_cast_1235_Sample/$exit
      -- CP-element group 459: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/type_cast_1235_sample_completed_
      -- 
    ra_3198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 459_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1235_inst_ack_0, ack => convTranspose_CP_39_elements(459)); -- 
    -- CP-element group 460:  transition  input  output  bypass 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	456 
    -- CP-element group 460: successors 
    -- CP-element group 460: 	461 
    -- CP-element group 460:  members (6) 
      -- CP-element group 460: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/type_cast_1235_Update/$exit
      -- CP-element group 460: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/type_cast_1235_Update/ca
      -- CP-element group 460: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/type_cast_1235_update_completed_
      -- CP-element group 460: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/WPIPE_elapsed_time_pipe_1242_Sample/req
      -- CP-element group 460: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/WPIPE_elapsed_time_pipe_1242_Sample/$entry
      -- CP-element group 460: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/WPIPE_elapsed_time_pipe_1242_sample_start_
      -- 
    ca_3203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 460_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1235_inst_ack_1, ack => convTranspose_CP_39_elements(460)); -- 
    req_3211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(460), ack => WPIPE_elapsed_time_pipe_1242_inst_req_0); -- 
    -- CP-element group 461:  transition  input  output  bypass 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	460 
    -- CP-element group 461: successors 
    -- CP-element group 461: 	462 
    -- CP-element group 461:  members (6) 
      -- CP-element group 461: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/WPIPE_elapsed_time_pipe_1242_Update/req
      -- CP-element group 461: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/WPIPE_elapsed_time_pipe_1242_Update/$entry
      -- CP-element group 461: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/WPIPE_elapsed_time_pipe_1242_Sample/ack
      -- CP-element group 461: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/WPIPE_elapsed_time_pipe_1242_Sample/$exit
      -- CP-element group 461: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/WPIPE_elapsed_time_pipe_1242_update_start_
      -- CP-element group 461: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/WPIPE_elapsed_time_pipe_1242_sample_completed_
      -- 
    ack_3212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 461_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1242_inst_ack_0, ack => convTranspose_CP_39_elements(461)); -- 
    req_3216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(461), ack => WPIPE_elapsed_time_pipe_1242_inst_req_1); -- 
    -- CP-element group 462:  branch  transition  place  input  output  bypass 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	461 
    -- CP-element group 462: successors 
    -- CP-element group 462: 	463 
    -- CP-element group 462: 	464 
    -- CP-element group 462:  members (13) 
      -- CP-element group 462: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244__exit__
      -- CP-element group 462: 	 branch_block_stmt_33/if_stmt_1246__entry__
      -- CP-element group 462: 	 branch_block_stmt_33/R_cmp408567_1247_place
      -- CP-element group 462: 	 branch_block_stmt_33/if_stmt_1246_else_link/$entry
      -- CP-element group 462: 	 branch_block_stmt_33/if_stmt_1246_if_link/$entry
      -- CP-element group 462: 	 branch_block_stmt_33/if_stmt_1246_eval_test/branch_req
      -- CP-element group 462: 	 branch_block_stmt_33/if_stmt_1246_eval_test/$exit
      -- CP-element group 462: 	 branch_block_stmt_33/if_stmt_1246_eval_test/$entry
      -- CP-element group 462: 	 branch_block_stmt_33/if_stmt_1246_dead_link/$entry
      -- CP-element group 462: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/WPIPE_elapsed_time_pipe_1242_Update/ack
      -- CP-element group 462: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/WPIPE_elapsed_time_pipe_1242_Update/$exit
      -- CP-element group 462: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/WPIPE_elapsed_time_pipe_1242_update_completed_
      -- CP-element group 462: 	 branch_block_stmt_33/call_stmt_1231_to_assign_stmt_1244/$exit
      -- 
    ack_3217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 462_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1242_inst_ack_1, ack => convTranspose_CP_39_elements(462)); -- 
    branch_req_3225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(462), ack => if_stmt_1246_branch_req_0); -- 
    -- CP-element group 463:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	462 
    -- CP-element group 463: successors 
    -- CP-element group 463: 	465 
    -- CP-element group 463: 	466 
    -- CP-element group 463:  members (18) 
      -- CP-element group 463: 	 branch_block_stmt_33/merge_stmt_1252__exit__
      -- CP-element group 463: 	 branch_block_stmt_33/assign_stmt_1258_to_assign_stmt_1287__entry__
      -- CP-element group 463: 	 branch_block_stmt_33/forx_xend417_bbx_xnph
      -- CP-element group 463: 	 branch_block_stmt_33/assign_stmt_1258_to_assign_stmt_1287/type_cast_1273_Update/cr
      -- CP-element group 463: 	 branch_block_stmt_33/assign_stmt_1258_to_assign_stmt_1287/type_cast_1273_Update/$entry
      -- CP-element group 463: 	 branch_block_stmt_33/assign_stmt_1258_to_assign_stmt_1287/type_cast_1273_Sample/rr
      -- CP-element group 463: 	 branch_block_stmt_33/assign_stmt_1258_to_assign_stmt_1287/type_cast_1273_Sample/$entry
      -- CP-element group 463: 	 branch_block_stmt_33/assign_stmt_1258_to_assign_stmt_1287/type_cast_1273_update_start_
      -- CP-element group 463: 	 branch_block_stmt_33/assign_stmt_1258_to_assign_stmt_1287/type_cast_1273_sample_start_
      -- CP-element group 463: 	 branch_block_stmt_33/assign_stmt_1258_to_assign_stmt_1287/$entry
      -- CP-element group 463: 	 branch_block_stmt_33/if_stmt_1246_if_link/if_choice_transition
      -- CP-element group 463: 	 branch_block_stmt_33/if_stmt_1246_if_link/$exit
      -- CP-element group 463: 	 branch_block_stmt_33/forx_xend417_bbx_xnph_PhiReq/$entry
      -- CP-element group 463: 	 branch_block_stmt_33/forx_xend417_bbx_xnph_PhiReq/$exit
      -- CP-element group 463: 	 branch_block_stmt_33/merge_stmt_1252_PhiReqMerge
      -- CP-element group 463: 	 branch_block_stmt_33/merge_stmt_1252_PhiAck/$entry
      -- CP-element group 463: 	 branch_block_stmt_33/merge_stmt_1252_PhiAck/$exit
      -- CP-element group 463: 	 branch_block_stmt_33/merge_stmt_1252_PhiAck/dummy
      -- 
    if_choice_transition_3230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 463_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1246_branch_ack_1, ack => convTranspose_CP_39_elements(463)); -- 
    cr_3252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(463), ack => type_cast_1273_inst_req_1); -- 
    rr_3247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(463), ack => type_cast_1273_inst_req_0); -- 
    -- CP-element group 464:  transition  place  input  bypass 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	462 
    -- CP-element group 464: successors 
    -- CP-element group 464: 	542 
    -- CP-element group 464:  members (5) 
      -- CP-element group 464: 	 branch_block_stmt_33/forx_xend417_forx_xend562
      -- CP-element group 464: 	 branch_block_stmt_33/if_stmt_1246_else_link/else_choice_transition
      -- CP-element group 464: 	 branch_block_stmt_33/if_stmt_1246_else_link/$exit
      -- CP-element group 464: 	 branch_block_stmt_33/forx_xend417_forx_xend562_PhiReq/$entry
      -- CP-element group 464: 	 branch_block_stmt_33/forx_xend417_forx_xend562_PhiReq/$exit
      -- 
    else_choice_transition_3234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 464_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1246_branch_ack_0, ack => convTranspose_CP_39_elements(464)); -- 
    -- CP-element group 465:  transition  input  bypass 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	463 
    -- CP-element group 465: successors 
    -- CP-element group 465:  members (3) 
      -- CP-element group 465: 	 branch_block_stmt_33/assign_stmt_1258_to_assign_stmt_1287/type_cast_1273_Sample/ra
      -- CP-element group 465: 	 branch_block_stmt_33/assign_stmt_1258_to_assign_stmt_1287/type_cast_1273_Sample/$exit
      -- CP-element group 465: 	 branch_block_stmt_33/assign_stmt_1258_to_assign_stmt_1287/type_cast_1273_sample_completed_
      -- 
    ra_3248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 465_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1273_inst_ack_0, ack => convTranspose_CP_39_elements(465)); -- 
    -- CP-element group 466:  transition  place  input  bypass 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	463 
    -- CP-element group 466: successors 
    -- CP-element group 466: 	536 
    -- CP-element group 466:  members (9) 
      -- CP-element group 466: 	 branch_block_stmt_33/assign_stmt_1258_to_assign_stmt_1287/type_cast_1273_Update/$exit
      -- CP-element group 466: 	 branch_block_stmt_33/assign_stmt_1258_to_assign_stmt_1287__exit__
      -- CP-element group 466: 	 branch_block_stmt_33/bbx_xnph_forx_xbody490
      -- CP-element group 466: 	 branch_block_stmt_33/assign_stmt_1258_to_assign_stmt_1287/type_cast_1273_Update/ca
      -- CP-element group 466: 	 branch_block_stmt_33/assign_stmt_1258_to_assign_stmt_1287/type_cast_1273_update_completed_
      -- CP-element group 466: 	 branch_block_stmt_33/assign_stmt_1258_to_assign_stmt_1287/$exit
      -- CP-element group 466: 	 branch_block_stmt_33/bbx_xnph_forx_xbody490_PhiReq/$entry
      -- CP-element group 466: 	 branch_block_stmt_33/bbx_xnph_forx_xbody490_PhiReq/phi_stmt_1290/$entry
      -- CP-element group 466: 	 branch_block_stmt_33/bbx_xnph_forx_xbody490_PhiReq/phi_stmt_1290/phi_stmt_1290_sources/$entry
      -- 
    ca_3253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 466_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1273_inst_ack_1, ack => convTranspose_CP_39_elements(466)); -- 
    -- CP-element group 467:  transition  input  bypass 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	541 
    -- CP-element group 467: successors 
    -- CP-element group 467: 	512 
    -- CP-element group 467:  members (3) 
      -- CP-element group 467: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_final_index_sum_regn_Sample/ack
      -- CP-element group 467: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_final_index_sum_regn_Sample/$exit
      -- CP-element group 467: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_final_index_sum_regn_sample_complete
      -- 
    ack_3282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 467_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1302_index_offset_ack_0, ack => convTranspose_CP_39_elements(467)); -- 
    -- CP-element group 468:  transition  input  output  bypass 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: 	541 
    -- CP-element group 468: successors 
    -- CP-element group 468: 	469 
    -- CP-element group 468:  members (11) 
      -- CP-element group 468: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_offset_calculated
      -- CP-element group 468: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_final_index_sum_regn_Update/ack
      -- CP-element group 468: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_base_plus_offset/sum_rename_req
      -- CP-element group 468: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/addr_of_1303_request/req
      -- CP-element group 468: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/addr_of_1303_sample_start_
      -- CP-element group 468: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_root_address_calculated
      -- CP-element group 468: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_base_plus_offset/sum_rename_ack
      -- CP-element group 468: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_final_index_sum_regn_Update/$exit
      -- CP-element group 468: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_base_plus_offset/$entry
      -- CP-element group 468: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_base_plus_offset/$exit
      -- CP-element group 468: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/addr_of_1303_request/$entry
      -- 
    ack_3287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 468_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1302_index_offset_ack_1, ack => convTranspose_CP_39_elements(468)); -- 
    req_3296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(468), ack => addr_of_1303_final_reg_req_0); -- 
    -- CP-element group 469:  transition  input  bypass 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	468 
    -- CP-element group 469: successors 
    -- CP-element group 469:  members (3) 
      -- CP-element group 469: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/addr_of_1303_request/ack
      -- CP-element group 469: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/addr_of_1303_sample_completed_
      -- CP-element group 469: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/addr_of_1303_request/$exit
      -- 
    ack_3297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 469_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1303_final_reg_ack_0, ack => convTranspose_CP_39_elements(469)); -- 
    -- CP-element group 470:  join  fork  transition  input  output  bypass 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	541 
    -- CP-element group 470: successors 
    -- CP-element group 470: 	471 
    -- CP-element group 470:  members (24) 
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_base_addr_resize/base_resize_req
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_base_plus_offset/sum_rename_req
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/addr_of_1303_update_completed_
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_base_addr_resize/$entry
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_base_addr_resize/$exit
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_base_address_calculated
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_word_address_calculated
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/addr_of_1303_complete/$exit
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_root_address_calculated
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/addr_of_1303_complete/ack
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_sample_start_
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_base_address_resized
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_base_addr_resize/base_resize_ack
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_base_plus_offset/$exit
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_base_plus_offset/$entry
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_Sample/word_access_start/word_0/rr
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_Sample/word_access_start/word_0/$entry
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_Sample/word_access_start/$entry
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_Sample/$entry
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_word_addrgen/root_register_ack
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_word_addrgen/root_register_req
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_word_addrgen/$exit
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_word_addrgen/$entry
      -- CP-element group 470: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_base_plus_offset/sum_rename_ack
      -- 
    ack_3302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 470_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1303_final_reg_ack_1, ack => convTranspose_CP_39_elements(470)); -- 
    rr_3335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(470), ack => ptr_deref_1307_load_0_req_0); -- 
    -- CP-element group 471:  transition  input  bypass 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	470 
    -- CP-element group 471: successors 
    -- CP-element group 471:  members (5) 
      -- CP-element group 471: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_sample_completed_
      -- CP-element group 471: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_Sample/word_access_start/word_0/ra
      -- CP-element group 471: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_Sample/word_access_start/word_0/$exit
      -- CP-element group 471: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_Sample/word_access_start/$exit
      -- CP-element group 471: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_Sample/$exit
      -- 
    ra_3336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 471_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1307_load_0_ack_0, ack => convTranspose_CP_39_elements(471)); -- 
    -- CP-element group 472:  fork  transition  input  output  bypass 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: 	541 
    -- CP-element group 472: successors 
    -- CP-element group 472: 	473 
    -- CP-element group 472: 	475 
    -- CP-element group 472: 	477 
    -- CP-element group 472: 	479 
    -- CP-element group 472: 	481 
    -- CP-element group 472: 	483 
    -- CP-element group 472: 	485 
    -- CP-element group 472: 	487 
    -- CP-element group 472:  members (33) 
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_update_completed_
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_Update/ptr_deref_1307_Merge/merge_ack
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_Update/ptr_deref_1307_Merge/merge_req
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_Update/ptr_deref_1307_Merge/$exit
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_Update/ptr_deref_1307_Merge/$entry
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_Update/word_access_complete/word_0/ca
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1311_sample_start_
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_Update/word_access_complete/word_0/$exit
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_Update/word_access_complete/$exit
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_Update/$exit
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1311_Sample/$entry
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1311_Sample/rr
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1321_sample_start_
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1321_Sample/$entry
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1321_Sample/rr
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1331_sample_start_
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1331_Sample/$entry
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1331_Sample/rr
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1341_sample_start_
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1341_Sample/$entry
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1341_Sample/rr
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1351_sample_start_
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1351_Sample/$entry
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1351_Sample/rr
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1361_sample_start_
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1361_Sample/$entry
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1361_Sample/rr
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1371_sample_start_
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1371_Sample/$entry
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1371_Sample/rr
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1381_sample_start_
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1381_Sample/$entry
      -- CP-element group 472: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1381_Sample/rr
      -- 
    ca_3347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 472_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1307_load_0_ack_1, ack => convTranspose_CP_39_elements(472)); -- 
    rr_3360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(472), ack => type_cast_1311_inst_req_0); -- 
    rr_3374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(472), ack => type_cast_1321_inst_req_0); -- 
    rr_3388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(472), ack => type_cast_1331_inst_req_0); -- 
    rr_3402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(472), ack => type_cast_1341_inst_req_0); -- 
    rr_3416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(472), ack => type_cast_1351_inst_req_0); -- 
    rr_3430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(472), ack => type_cast_1361_inst_req_0); -- 
    rr_3444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(472), ack => type_cast_1371_inst_req_0); -- 
    rr_3458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(472), ack => type_cast_1381_inst_req_0); -- 
    -- CP-element group 473:  transition  input  bypass 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	472 
    -- CP-element group 473: successors 
    -- CP-element group 473:  members (3) 
      -- CP-element group 473: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1311_sample_completed_
      -- CP-element group 473: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1311_Sample/$exit
      -- CP-element group 473: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1311_Sample/ra
      -- 
    ra_3361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 473_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1311_inst_ack_0, ack => convTranspose_CP_39_elements(473)); -- 
    -- CP-element group 474:  transition  input  bypass 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	541 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	509 
    -- CP-element group 474:  members (3) 
      -- CP-element group 474: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1311_update_completed_
      -- CP-element group 474: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1311_Update/$exit
      -- CP-element group 474: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1311_Update/ca
      -- 
    ca_3366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 474_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1311_inst_ack_1, ack => convTranspose_CP_39_elements(474)); -- 
    -- CP-element group 475:  transition  input  bypass 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	472 
    -- CP-element group 475: successors 
    -- CP-element group 475:  members (3) 
      -- CP-element group 475: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1321_sample_completed_
      -- CP-element group 475: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1321_Sample/$exit
      -- CP-element group 475: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1321_Sample/ra
      -- 
    ra_3375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 475_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1321_inst_ack_0, ack => convTranspose_CP_39_elements(475)); -- 
    -- CP-element group 476:  transition  input  bypass 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: 	541 
    -- CP-element group 476: successors 
    -- CP-element group 476: 	506 
    -- CP-element group 476:  members (3) 
      -- CP-element group 476: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1321_update_completed_
      -- CP-element group 476: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1321_Update/$exit
      -- CP-element group 476: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1321_Update/ca
      -- 
    ca_3380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 476_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1321_inst_ack_1, ack => convTranspose_CP_39_elements(476)); -- 
    -- CP-element group 477:  transition  input  bypass 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	472 
    -- CP-element group 477: successors 
    -- CP-element group 477:  members (3) 
      -- CP-element group 477: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1331_sample_completed_
      -- CP-element group 477: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1331_Sample/$exit
      -- CP-element group 477: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1331_Sample/ra
      -- 
    ra_3389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 477_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1331_inst_ack_0, ack => convTranspose_CP_39_elements(477)); -- 
    -- CP-element group 478:  transition  input  bypass 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: 	541 
    -- CP-element group 478: successors 
    -- CP-element group 478: 	503 
    -- CP-element group 478:  members (3) 
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1331_update_completed_
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1331_Update/$exit
      -- CP-element group 478: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1331_Update/ca
      -- 
    ca_3394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 478_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1331_inst_ack_1, ack => convTranspose_CP_39_elements(478)); -- 
    -- CP-element group 479:  transition  input  bypass 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	472 
    -- CP-element group 479: successors 
    -- CP-element group 479:  members (3) 
      -- CP-element group 479: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1341_sample_completed_
      -- CP-element group 479: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1341_Sample/$exit
      -- CP-element group 479: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1341_Sample/ra
      -- 
    ra_3403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 479_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1341_inst_ack_0, ack => convTranspose_CP_39_elements(479)); -- 
    -- CP-element group 480:  transition  input  bypass 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: 	541 
    -- CP-element group 480: successors 
    -- CP-element group 480: 	500 
    -- CP-element group 480:  members (3) 
      -- CP-element group 480: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1341_update_completed_
      -- CP-element group 480: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1341_Update/$exit
      -- CP-element group 480: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1341_Update/ca
      -- 
    ca_3408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 480_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1341_inst_ack_1, ack => convTranspose_CP_39_elements(480)); -- 
    -- CP-element group 481:  transition  input  bypass 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	472 
    -- CP-element group 481: successors 
    -- CP-element group 481:  members (3) 
      -- CP-element group 481: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1351_sample_completed_
      -- CP-element group 481: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1351_Sample/$exit
      -- CP-element group 481: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1351_Sample/ra
      -- 
    ra_3417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 481_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1351_inst_ack_0, ack => convTranspose_CP_39_elements(481)); -- 
    -- CP-element group 482:  transition  input  bypass 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	541 
    -- CP-element group 482: successors 
    -- CP-element group 482: 	497 
    -- CP-element group 482:  members (3) 
      -- CP-element group 482: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1351_update_completed_
      -- CP-element group 482: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1351_Update/$exit
      -- CP-element group 482: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1351_Update/ca
      -- 
    ca_3422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 482_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1351_inst_ack_1, ack => convTranspose_CP_39_elements(482)); -- 
    -- CP-element group 483:  transition  input  bypass 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: 	472 
    -- CP-element group 483: successors 
    -- CP-element group 483:  members (3) 
      -- CP-element group 483: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1361_sample_completed_
      -- CP-element group 483: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1361_Sample/$exit
      -- CP-element group 483: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1361_Sample/ra
      -- 
    ra_3431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 483_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1361_inst_ack_0, ack => convTranspose_CP_39_elements(483)); -- 
    -- CP-element group 484:  transition  input  bypass 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	541 
    -- CP-element group 484: successors 
    -- CP-element group 484: 	494 
    -- CP-element group 484:  members (3) 
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1361_update_completed_
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1361_Update/$exit
      -- CP-element group 484: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1361_Update/ca
      -- 
    ca_3436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 484_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1361_inst_ack_1, ack => convTranspose_CP_39_elements(484)); -- 
    -- CP-element group 485:  transition  input  bypass 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	472 
    -- CP-element group 485: successors 
    -- CP-element group 485:  members (3) 
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1371_sample_completed_
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1371_Sample/$exit
      -- CP-element group 485: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1371_Sample/ra
      -- 
    ra_3445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 485_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1371_inst_ack_0, ack => convTranspose_CP_39_elements(485)); -- 
    -- CP-element group 486:  transition  input  bypass 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: 	541 
    -- CP-element group 486: successors 
    -- CP-element group 486: 	491 
    -- CP-element group 486:  members (3) 
      -- CP-element group 486: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1371_update_completed_
      -- CP-element group 486: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1371_Update/$exit
      -- CP-element group 486: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1371_Update/ca
      -- 
    ca_3450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 486_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1371_inst_ack_1, ack => convTranspose_CP_39_elements(486)); -- 
    -- CP-element group 487:  transition  input  bypass 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: 	472 
    -- CP-element group 487: successors 
    -- CP-element group 487:  members (3) 
      -- CP-element group 487: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1381_sample_completed_
      -- CP-element group 487: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1381_Sample/$exit
      -- CP-element group 487: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1381_Sample/ra
      -- 
    ra_3459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 487_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1381_inst_ack_0, ack => convTranspose_CP_39_elements(487)); -- 
    -- CP-element group 488:  transition  input  output  bypass 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: 	541 
    -- CP-element group 488: successors 
    -- CP-element group 488: 	489 
    -- CP-element group 488:  members (6) 
      -- CP-element group 488: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1381_update_completed_
      -- CP-element group 488: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1381_Update/$exit
      -- CP-element group 488: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1381_Update/ca
      -- CP-element group 488: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1383_sample_start_
      -- CP-element group 488: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1383_Sample/$entry
      -- CP-element group 488: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1383_Sample/req
      -- 
    ca_3464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 488_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1381_inst_ack_1, ack => convTranspose_CP_39_elements(488)); -- 
    req_3472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(488), ack => WPIPE_ConvTranspose_output_pipe_1383_inst_req_0); -- 
    -- CP-element group 489:  transition  input  output  bypass 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	488 
    -- CP-element group 489: successors 
    -- CP-element group 489: 	490 
    -- CP-element group 489:  members (6) 
      -- CP-element group 489: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1383_sample_completed_
      -- CP-element group 489: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1383_update_start_
      -- CP-element group 489: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1383_Sample/$exit
      -- CP-element group 489: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1383_Sample/ack
      -- CP-element group 489: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1383_Update/$entry
      -- CP-element group 489: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1383_Update/req
      -- 
    ack_3473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 489_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1383_inst_ack_0, ack => convTranspose_CP_39_elements(489)); -- 
    req_3477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => WPIPE_ConvTranspose_output_pipe_1383_inst_req_1); -- 
    -- CP-element group 490:  transition  input  bypass 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: 	489 
    -- CP-element group 490: successors 
    -- CP-element group 490: 	491 
    -- CP-element group 490:  members (3) 
      -- CP-element group 490: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1383_update_completed_
      -- CP-element group 490: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1383_Update/$exit
      -- CP-element group 490: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1383_Update/ack
      -- 
    ack_3478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 490_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1383_inst_ack_1, ack => convTranspose_CP_39_elements(490)); -- 
    -- CP-element group 491:  join  transition  output  bypass 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: 	486 
    -- CP-element group 491: 	490 
    -- CP-element group 491: successors 
    -- CP-element group 491: 	492 
    -- CP-element group 491:  members (3) 
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1386_sample_start_
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1386_Sample/$entry
      -- CP-element group 491: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1386_Sample/req
      -- 
    req_3486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(491), ack => WPIPE_ConvTranspose_output_pipe_1386_inst_req_0); -- 
    convTranspose_cp_element_group_491: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_491"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(486) & convTranspose_CP_39_elements(490);
      gj_convTranspose_cp_element_group_491 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(491), clk => clk, reset => reset); --
    end block;
    -- CP-element group 492:  transition  input  output  bypass 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: 	491 
    -- CP-element group 492: successors 
    -- CP-element group 492: 	493 
    -- CP-element group 492:  members (6) 
      -- CP-element group 492: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1386_sample_completed_
      -- CP-element group 492: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1386_update_start_
      -- CP-element group 492: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1386_Sample/$exit
      -- CP-element group 492: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1386_Sample/ack
      -- CP-element group 492: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1386_Update/$entry
      -- CP-element group 492: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1386_Update/req
      -- 
    ack_3487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 492_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1386_inst_ack_0, ack => convTranspose_CP_39_elements(492)); -- 
    req_3491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(492), ack => WPIPE_ConvTranspose_output_pipe_1386_inst_req_1); -- 
    -- CP-element group 493:  transition  input  bypass 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	492 
    -- CP-element group 493: successors 
    -- CP-element group 493: 	494 
    -- CP-element group 493:  members (3) 
      -- CP-element group 493: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1386_update_completed_
      -- CP-element group 493: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1386_Update/$exit
      -- CP-element group 493: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1386_Update/ack
      -- 
    ack_3492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 493_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1386_inst_ack_1, ack => convTranspose_CP_39_elements(493)); -- 
    -- CP-element group 494:  join  transition  output  bypass 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	493 
    -- CP-element group 494: 	484 
    -- CP-element group 494: successors 
    -- CP-element group 494: 	495 
    -- CP-element group 494:  members (3) 
      -- CP-element group 494: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1389_sample_start_
      -- CP-element group 494: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1389_Sample/$entry
      -- CP-element group 494: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1389_Sample/req
      -- 
    req_3500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(494), ack => WPIPE_ConvTranspose_output_pipe_1389_inst_req_0); -- 
    convTranspose_cp_element_group_494: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_494"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(493) & convTranspose_CP_39_elements(484);
      gj_convTranspose_cp_element_group_494 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(494), clk => clk, reset => reset); --
    end block;
    -- CP-element group 495:  transition  input  output  bypass 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	494 
    -- CP-element group 495: successors 
    -- CP-element group 495: 	496 
    -- CP-element group 495:  members (6) 
      -- CP-element group 495: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1389_sample_completed_
      -- CP-element group 495: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1389_update_start_
      -- CP-element group 495: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1389_Sample/$exit
      -- CP-element group 495: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1389_Sample/ack
      -- CP-element group 495: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1389_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1389_Update/req
      -- 
    ack_3501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 495_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1389_inst_ack_0, ack => convTranspose_CP_39_elements(495)); -- 
    req_3505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => WPIPE_ConvTranspose_output_pipe_1389_inst_req_1); -- 
    -- CP-element group 496:  transition  input  bypass 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	495 
    -- CP-element group 496: successors 
    -- CP-element group 496: 	497 
    -- CP-element group 496:  members (3) 
      -- CP-element group 496: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1389_update_completed_
      -- CP-element group 496: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1389_Update/$exit
      -- CP-element group 496: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1389_Update/ack
      -- 
    ack_3506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 496_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1389_inst_ack_1, ack => convTranspose_CP_39_elements(496)); -- 
    -- CP-element group 497:  join  transition  output  bypass 
    -- CP-element group 497: predecessors 
    -- CP-element group 497: 	496 
    -- CP-element group 497: 	482 
    -- CP-element group 497: successors 
    -- CP-element group 497: 	498 
    -- CP-element group 497:  members (3) 
      -- CP-element group 497: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1392_sample_start_
      -- CP-element group 497: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1392_Sample/$entry
      -- CP-element group 497: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1392_Sample/req
      -- 
    req_3514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(497), ack => WPIPE_ConvTranspose_output_pipe_1392_inst_req_0); -- 
    convTranspose_cp_element_group_497: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_497"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(496) & convTranspose_CP_39_elements(482);
      gj_convTranspose_cp_element_group_497 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(497), clk => clk, reset => reset); --
    end block;
    -- CP-element group 498:  transition  input  output  bypass 
    -- CP-element group 498: predecessors 
    -- CP-element group 498: 	497 
    -- CP-element group 498: successors 
    -- CP-element group 498: 	499 
    -- CP-element group 498:  members (6) 
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1392_sample_completed_
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1392_update_start_
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1392_Sample/$exit
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1392_Sample/ack
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1392_Update/$entry
      -- CP-element group 498: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1392_Update/req
      -- 
    ack_3515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 498_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1392_inst_ack_0, ack => convTranspose_CP_39_elements(498)); -- 
    req_3519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(498), ack => WPIPE_ConvTranspose_output_pipe_1392_inst_req_1); -- 
    -- CP-element group 499:  transition  input  bypass 
    -- CP-element group 499: predecessors 
    -- CP-element group 499: 	498 
    -- CP-element group 499: successors 
    -- CP-element group 499: 	500 
    -- CP-element group 499:  members (3) 
      -- CP-element group 499: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1392_update_completed_
      -- CP-element group 499: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1392_Update/$exit
      -- CP-element group 499: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1392_Update/ack
      -- 
    ack_3520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 499_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1392_inst_ack_1, ack => convTranspose_CP_39_elements(499)); -- 
    -- CP-element group 500:  join  transition  output  bypass 
    -- CP-element group 500: predecessors 
    -- CP-element group 500: 	499 
    -- CP-element group 500: 	480 
    -- CP-element group 500: successors 
    -- CP-element group 500: 	501 
    -- CP-element group 500:  members (3) 
      -- CP-element group 500: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1395_sample_start_
      -- CP-element group 500: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1395_Sample/$entry
      -- CP-element group 500: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1395_Sample/req
      -- 
    req_3528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(500), ack => WPIPE_ConvTranspose_output_pipe_1395_inst_req_0); -- 
    convTranspose_cp_element_group_500: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_500"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(499) & convTranspose_CP_39_elements(480);
      gj_convTranspose_cp_element_group_500 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(500), clk => clk, reset => reset); --
    end block;
    -- CP-element group 501:  transition  input  output  bypass 
    -- CP-element group 501: predecessors 
    -- CP-element group 501: 	500 
    -- CP-element group 501: successors 
    -- CP-element group 501: 	502 
    -- CP-element group 501:  members (6) 
      -- CP-element group 501: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1395_sample_completed_
      -- CP-element group 501: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1395_update_start_
      -- CP-element group 501: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1395_Sample/$exit
      -- CP-element group 501: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1395_Sample/ack
      -- CP-element group 501: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1395_Update/$entry
      -- CP-element group 501: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1395_Update/req
      -- 
    ack_3529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 501_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1395_inst_ack_0, ack => convTranspose_CP_39_elements(501)); -- 
    req_3533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(501), ack => WPIPE_ConvTranspose_output_pipe_1395_inst_req_1); -- 
    -- CP-element group 502:  transition  input  bypass 
    -- CP-element group 502: predecessors 
    -- CP-element group 502: 	501 
    -- CP-element group 502: successors 
    -- CP-element group 502: 	503 
    -- CP-element group 502:  members (3) 
      -- CP-element group 502: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1395_update_completed_
      -- CP-element group 502: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1395_Update/$exit
      -- CP-element group 502: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1395_Update/ack
      -- 
    ack_3534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 502_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1395_inst_ack_1, ack => convTranspose_CP_39_elements(502)); -- 
    -- CP-element group 503:  join  transition  output  bypass 
    -- CP-element group 503: predecessors 
    -- CP-element group 503: 	502 
    -- CP-element group 503: 	478 
    -- CP-element group 503: successors 
    -- CP-element group 503: 	504 
    -- CP-element group 503:  members (3) 
      -- CP-element group 503: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1398_sample_start_
      -- CP-element group 503: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1398_Sample/$entry
      -- CP-element group 503: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1398_Sample/req
      -- 
    req_3542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(503), ack => WPIPE_ConvTranspose_output_pipe_1398_inst_req_0); -- 
    convTranspose_cp_element_group_503: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_503"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(502) & convTranspose_CP_39_elements(478);
      gj_convTranspose_cp_element_group_503 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(503), clk => clk, reset => reset); --
    end block;
    -- CP-element group 504:  transition  input  output  bypass 
    -- CP-element group 504: predecessors 
    -- CP-element group 504: 	503 
    -- CP-element group 504: successors 
    -- CP-element group 504: 	505 
    -- CP-element group 504:  members (6) 
      -- CP-element group 504: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1398_sample_completed_
      -- CP-element group 504: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1398_update_start_
      -- CP-element group 504: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1398_Sample/$exit
      -- CP-element group 504: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1398_Sample/ack
      -- CP-element group 504: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1398_Update/$entry
      -- CP-element group 504: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1398_Update/req
      -- 
    ack_3543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 504_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1398_inst_ack_0, ack => convTranspose_CP_39_elements(504)); -- 
    req_3547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(504), ack => WPIPE_ConvTranspose_output_pipe_1398_inst_req_1); -- 
    -- CP-element group 505:  transition  input  bypass 
    -- CP-element group 505: predecessors 
    -- CP-element group 505: 	504 
    -- CP-element group 505: successors 
    -- CP-element group 505: 	506 
    -- CP-element group 505:  members (3) 
      -- CP-element group 505: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1398_update_completed_
      -- CP-element group 505: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1398_Update/$exit
      -- CP-element group 505: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1398_Update/ack
      -- 
    ack_3548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 505_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1398_inst_ack_1, ack => convTranspose_CP_39_elements(505)); -- 
    -- CP-element group 506:  join  transition  output  bypass 
    -- CP-element group 506: predecessors 
    -- CP-element group 506: 	505 
    -- CP-element group 506: 	476 
    -- CP-element group 506: successors 
    -- CP-element group 506: 	507 
    -- CP-element group 506:  members (3) 
      -- CP-element group 506: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1401_sample_start_
      -- CP-element group 506: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1401_Sample/$entry
      -- CP-element group 506: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1401_Sample/req
      -- 
    req_3556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(506), ack => WPIPE_ConvTranspose_output_pipe_1401_inst_req_0); -- 
    convTranspose_cp_element_group_506: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_506"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(505) & convTranspose_CP_39_elements(476);
      gj_convTranspose_cp_element_group_506 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(506), clk => clk, reset => reset); --
    end block;
    -- CP-element group 507:  transition  input  output  bypass 
    -- CP-element group 507: predecessors 
    -- CP-element group 507: 	506 
    -- CP-element group 507: successors 
    -- CP-element group 507: 	508 
    -- CP-element group 507:  members (6) 
      -- CP-element group 507: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1401_sample_completed_
      -- CP-element group 507: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1401_update_start_
      -- CP-element group 507: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1401_Sample/$exit
      -- CP-element group 507: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1401_Sample/ack
      -- CP-element group 507: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1401_Update/$entry
      -- CP-element group 507: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1401_Update/req
      -- 
    ack_3557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 507_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1401_inst_ack_0, ack => convTranspose_CP_39_elements(507)); -- 
    req_3561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(507), ack => WPIPE_ConvTranspose_output_pipe_1401_inst_req_1); -- 
    -- CP-element group 508:  transition  input  bypass 
    -- CP-element group 508: predecessors 
    -- CP-element group 508: 	507 
    -- CP-element group 508: successors 
    -- CP-element group 508: 	509 
    -- CP-element group 508:  members (3) 
      -- CP-element group 508: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1401_update_completed_
      -- CP-element group 508: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1401_Update/$exit
      -- CP-element group 508: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1401_Update/ack
      -- 
    ack_3562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 508_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1401_inst_ack_1, ack => convTranspose_CP_39_elements(508)); -- 
    -- CP-element group 509:  join  transition  output  bypass 
    -- CP-element group 509: predecessors 
    -- CP-element group 509: 	508 
    -- CP-element group 509: 	474 
    -- CP-element group 509: successors 
    -- CP-element group 509: 	510 
    -- CP-element group 509:  members (3) 
      -- CP-element group 509: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1404_sample_start_
      -- CP-element group 509: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1404_Sample/$entry
      -- CP-element group 509: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1404_Sample/req
      -- 
    req_3570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(509), ack => WPIPE_ConvTranspose_output_pipe_1404_inst_req_0); -- 
    convTranspose_cp_element_group_509: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_509"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(508) & convTranspose_CP_39_elements(474);
      gj_convTranspose_cp_element_group_509 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(509), clk => clk, reset => reset); --
    end block;
    -- CP-element group 510:  transition  input  output  bypass 
    -- CP-element group 510: predecessors 
    -- CP-element group 510: 	509 
    -- CP-element group 510: successors 
    -- CP-element group 510: 	511 
    -- CP-element group 510:  members (6) 
      -- CP-element group 510: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1404_sample_completed_
      -- CP-element group 510: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1404_update_start_
      -- CP-element group 510: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1404_Sample/$exit
      -- CP-element group 510: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1404_Sample/ack
      -- CP-element group 510: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1404_Update/$entry
      -- CP-element group 510: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1404_Update/req
      -- 
    ack_3571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 510_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1404_inst_ack_0, ack => convTranspose_CP_39_elements(510)); -- 
    req_3575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(510), ack => WPIPE_ConvTranspose_output_pipe_1404_inst_req_1); -- 
    -- CP-element group 511:  transition  input  bypass 
    -- CP-element group 511: predecessors 
    -- CP-element group 511: 	510 
    -- CP-element group 511: successors 
    -- CP-element group 511: 	512 
    -- CP-element group 511:  members (3) 
      -- CP-element group 511: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1404_update_completed_
      -- CP-element group 511: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1404_Update/$exit
      -- CP-element group 511: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/WPIPE_ConvTranspose_output_pipe_1404_Update/ack
      -- 
    ack_3576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 511_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1404_inst_ack_1, ack => convTranspose_CP_39_elements(511)); -- 
    -- CP-element group 512:  branch  join  transition  place  output  bypass 
    -- CP-element group 512: predecessors 
    -- CP-element group 512: 	511 
    -- CP-element group 512: 	467 
    -- CP-element group 512: successors 
    -- CP-element group 512: 	513 
    -- CP-element group 512: 	514 
    -- CP-element group 512:  members (10) 
      -- CP-element group 512: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417__exit__
      -- CP-element group 512: 	 branch_block_stmt_33/if_stmt_1418__entry__
      -- CP-element group 512: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/$exit
      -- CP-element group 512: 	 branch_block_stmt_33/if_stmt_1418_dead_link/$entry
      -- CP-element group 512: 	 branch_block_stmt_33/if_stmt_1418_eval_test/$entry
      -- CP-element group 512: 	 branch_block_stmt_33/if_stmt_1418_eval_test/$exit
      -- CP-element group 512: 	 branch_block_stmt_33/if_stmt_1418_eval_test/branch_req
      -- CP-element group 512: 	 branch_block_stmt_33/R_exitcond1_1419_place
      -- CP-element group 512: 	 branch_block_stmt_33/if_stmt_1418_if_link/$entry
      -- CP-element group 512: 	 branch_block_stmt_33/if_stmt_1418_else_link/$entry
      -- 
    branch_req_3584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(512), ack => if_stmt_1418_branch_req_0); -- 
    convTranspose_cp_element_group_512: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_512"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(511) & convTranspose_CP_39_elements(467);
      gj_convTranspose_cp_element_group_512 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(512), clk => clk, reset => reset); --
    end block;
    -- CP-element group 513:  merge  transition  place  input  bypass 
    -- CP-element group 513: predecessors 
    -- CP-element group 513: 	512 
    -- CP-element group 513: successors 
    -- CP-element group 513: 	542 
    -- CP-element group 513:  members (13) 
      -- CP-element group 513: 	 branch_block_stmt_33/merge_stmt_1424__exit__
      -- CP-element group 513: 	 branch_block_stmt_33/forx_xend562x_xloopexit_forx_xend562
      -- CP-element group 513: 	 branch_block_stmt_33/if_stmt_1418_if_link/$exit
      -- CP-element group 513: 	 branch_block_stmt_33/if_stmt_1418_if_link/if_choice_transition
      -- CP-element group 513: 	 branch_block_stmt_33/forx_xbody490_forx_xend562x_xloopexit
      -- CP-element group 513: 	 branch_block_stmt_33/forx_xbody490_forx_xend562x_xloopexit_PhiReq/$entry
      -- CP-element group 513: 	 branch_block_stmt_33/forx_xbody490_forx_xend562x_xloopexit_PhiReq/$exit
      -- CP-element group 513: 	 branch_block_stmt_33/merge_stmt_1424_PhiReqMerge
      -- CP-element group 513: 	 branch_block_stmt_33/merge_stmt_1424_PhiAck/$entry
      -- CP-element group 513: 	 branch_block_stmt_33/merge_stmt_1424_PhiAck/$exit
      -- CP-element group 513: 	 branch_block_stmt_33/merge_stmt_1424_PhiAck/dummy
      -- CP-element group 513: 	 branch_block_stmt_33/forx_xend562x_xloopexit_forx_xend562_PhiReq/$entry
      -- CP-element group 513: 	 branch_block_stmt_33/forx_xend562x_xloopexit_forx_xend562_PhiReq/$exit
      -- 
    if_choice_transition_3589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 513_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1418_branch_ack_1, ack => convTranspose_CP_39_elements(513)); -- 
    -- CP-element group 514:  fork  transition  place  input  output  bypass 
    -- CP-element group 514: predecessors 
    -- CP-element group 514: 	512 
    -- CP-element group 514: successors 
    -- CP-element group 514: 	538 
    -- CP-element group 514: 	537 
    -- CP-element group 514:  members (12) 
      -- CP-element group 514: 	 branch_block_stmt_33/if_stmt_1418_else_link/$exit
      -- CP-element group 514: 	 branch_block_stmt_33/if_stmt_1418_else_link/else_choice_transition
      -- CP-element group 514: 	 branch_block_stmt_33/forx_xbody490_forx_xbody490
      -- CP-element group 514: 	 branch_block_stmt_33/forx_xbody490_forx_xbody490_PhiReq/$entry
      -- CP-element group 514: 	 branch_block_stmt_33/forx_xbody490_forx_xbody490_PhiReq/phi_stmt_1290/$entry
      -- CP-element group 514: 	 branch_block_stmt_33/forx_xbody490_forx_xbody490_PhiReq/phi_stmt_1290/phi_stmt_1290_sources/$entry
      -- CP-element group 514: 	 branch_block_stmt_33/forx_xbody490_forx_xbody490_PhiReq/phi_stmt_1290/phi_stmt_1290_sources/type_cast_1293/$entry
      -- CP-element group 514: 	 branch_block_stmt_33/forx_xbody490_forx_xbody490_PhiReq/phi_stmt_1290/phi_stmt_1290_sources/type_cast_1293/SplitProtocol/$entry
      -- CP-element group 514: 	 branch_block_stmt_33/forx_xbody490_forx_xbody490_PhiReq/phi_stmt_1290/phi_stmt_1290_sources/type_cast_1293/SplitProtocol/Sample/$entry
      -- CP-element group 514: 	 branch_block_stmt_33/forx_xbody490_forx_xbody490_PhiReq/phi_stmt_1290/phi_stmt_1290_sources/type_cast_1293/SplitProtocol/Sample/rr
      -- CP-element group 514: 	 branch_block_stmt_33/forx_xbody490_forx_xbody490_PhiReq/phi_stmt_1290/phi_stmt_1290_sources/type_cast_1293/SplitProtocol/Update/$entry
      -- CP-element group 514: 	 branch_block_stmt_33/forx_xbody490_forx_xbody490_PhiReq/phi_stmt_1290/phi_stmt_1290_sources/type_cast_1293/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 514_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1418_branch_ack_0, ack => convTranspose_CP_39_elements(514)); -- 
    rr_3868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(514), ack => type_cast_1293_inst_req_0); -- 
    cr_3873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(514), ack => type_cast_1293_inst_req_1); -- 
    -- CP-element group 515:  merge  branch  transition  place  output  bypass 
    -- CP-element group 515: predecessors 
    -- CP-element group 515: 	191 
    -- CP-element group 515: 	259 
    -- CP-element group 515: successors 
    -- CP-element group 515: 	192 
    -- CP-element group 515: 	193 
    -- CP-element group 515:  members (17) 
      -- CP-element group 515: 	 branch_block_stmt_33/merge_stmt_474__exit__
      -- CP-element group 515: 	 branch_block_stmt_33/assign_stmt_480__entry__
      -- CP-element group 515: 	 branch_block_stmt_33/assign_stmt_480__exit__
      -- CP-element group 515: 	 branch_block_stmt_33/if_stmt_481__entry__
      -- CP-element group 515: 	 branch_block_stmt_33/if_stmt_481_else_link/$entry
      -- CP-element group 515: 	 branch_block_stmt_33/if_stmt_481_if_link/$entry
      -- CP-element group 515: 	 branch_block_stmt_33/R_cmp306571_482_place
      -- CP-element group 515: 	 branch_block_stmt_33/if_stmt_481_eval_test/branch_req
      -- CP-element group 515: 	 branch_block_stmt_33/if_stmt_481_eval_test/$exit
      -- CP-element group 515: 	 branch_block_stmt_33/if_stmt_481_eval_test/$entry
      -- CP-element group 515: 	 branch_block_stmt_33/if_stmt_481_dead_link/$entry
      -- CP-element group 515: 	 branch_block_stmt_33/assign_stmt_480/$exit
      -- CP-element group 515: 	 branch_block_stmt_33/assign_stmt_480/$entry
      -- CP-element group 515: 	 branch_block_stmt_33/merge_stmt_474_PhiReqMerge
      -- CP-element group 515: 	 branch_block_stmt_33/merge_stmt_474_PhiAck/$entry
      -- CP-element group 515: 	 branch_block_stmt_33/merge_stmt_474_PhiAck/$exit
      -- CP-element group 515: 	 branch_block_stmt_33/merge_stmt_474_PhiAck/dummy
      -- 
    branch_req_1261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(515), ack => if_stmt_481_branch_req_0); -- 
    convTranspose_CP_39_elements(515) <= OrReduce(convTranspose_CP_39_elements(191) & convTranspose_CP_39_elements(259));
    -- CP-element group 516:  transition  output  delay-element  bypass 
    -- CP-element group 516: predecessors 
    -- CP-element group 516: 	195 
    -- CP-element group 516: successors 
    -- CP-element group 516: 	520 
    -- CP-element group 516:  members (5) 
      -- CP-element group 516: 	 branch_block_stmt_33/bbx_xnph577_forx_xbody_PhiReq/$exit
      -- CP-element group 516: 	 branch_block_stmt_33/bbx_xnph577_forx_xbody_PhiReq/phi_stmt_525/$exit
      -- CP-element group 516: 	 branch_block_stmt_33/bbx_xnph577_forx_xbody_PhiReq/phi_stmt_525/phi_stmt_525_sources/$exit
      -- CP-element group 516: 	 branch_block_stmt_33/bbx_xnph577_forx_xbody_PhiReq/phi_stmt_525/phi_stmt_525_sources/type_cast_529_konst_delay_trans
      -- CP-element group 516: 	 branch_block_stmt_33/bbx_xnph577_forx_xbody_PhiReq/phi_stmt_525/phi_stmt_525_req
      -- 
    phi_stmt_525_req_3641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_525_req_3641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(516), ack => phi_stmt_525_req_0); -- 
    -- Element group convTranspose_CP_39_elements(516) is a control-delay.
    cp_element_516_delay: control_delay_element  generic map(name => " 516_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(195), ack => convTranspose_CP_39_elements(516), clk => clk, reset =>reset);
    -- CP-element group 517:  transition  input  bypass 
    -- CP-element group 517: predecessors 
    -- CP-element group 517: 	260 
    -- CP-element group 517: successors 
    -- CP-element group 517: 	519 
    -- CP-element group 517:  members (2) 
      -- CP-element group 517: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_525/phi_stmt_525_sources/type_cast_531/SplitProtocol/Sample/$exit
      -- CP-element group 517: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_525/phi_stmt_525_sources/type_cast_531/SplitProtocol/Sample/ra
      -- 
    ra_3661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 517_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_531_inst_ack_0, ack => convTranspose_CP_39_elements(517)); -- 
    -- CP-element group 518:  transition  input  bypass 
    -- CP-element group 518: predecessors 
    -- CP-element group 518: 	260 
    -- CP-element group 518: successors 
    -- CP-element group 518: 	519 
    -- CP-element group 518:  members (2) 
      -- CP-element group 518: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_525/phi_stmt_525_sources/type_cast_531/SplitProtocol/Update/$exit
      -- CP-element group 518: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_525/phi_stmt_525_sources/type_cast_531/SplitProtocol/Update/ca
      -- 
    ca_3666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 518_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_531_inst_ack_1, ack => convTranspose_CP_39_elements(518)); -- 
    -- CP-element group 519:  join  transition  output  bypass 
    -- CP-element group 519: predecessors 
    -- CP-element group 519: 	517 
    -- CP-element group 519: 	518 
    -- CP-element group 519: successors 
    -- CP-element group 519: 	520 
    -- CP-element group 519:  members (6) 
      -- CP-element group 519: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 519: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_525/$exit
      -- CP-element group 519: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_525/phi_stmt_525_sources/$exit
      -- CP-element group 519: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_525/phi_stmt_525_sources/type_cast_531/$exit
      -- CP-element group 519: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_525/phi_stmt_525_sources/type_cast_531/SplitProtocol/$exit
      -- CP-element group 519: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_525/phi_stmt_525_req
      -- 
    phi_stmt_525_req_3667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_525_req_3667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(519), ack => phi_stmt_525_req_1); -- 
    convTranspose_cp_element_group_519: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_519"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(517) & convTranspose_CP_39_elements(518);
      gj_convTranspose_cp_element_group_519 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(519), clk => clk, reset => reset); --
    end block;
    -- CP-element group 520:  merge  transition  place  bypass 
    -- CP-element group 520: predecessors 
    -- CP-element group 520: 	516 
    -- CP-element group 520: 	519 
    -- CP-element group 520: successors 
    -- CP-element group 520: 	521 
    -- CP-element group 520:  members (2) 
      -- CP-element group 520: 	 branch_block_stmt_33/merge_stmt_524_PhiReqMerge
      -- CP-element group 520: 	 branch_block_stmt_33/merge_stmt_524_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(520) <= OrReduce(convTranspose_CP_39_elements(516) & convTranspose_CP_39_elements(519));
    -- CP-element group 521:  fork  transition  place  input  output  bypass 
    -- CP-element group 521: predecessors 
    -- CP-element group 521: 	520 
    -- CP-element group 521: successors 
    -- CP-element group 521: 	196 
    -- CP-element group 521: 	197 
    -- CP-element group 521: 	199 
    -- CP-element group 521: 	200 
    -- CP-element group 521: 	205 
    -- CP-element group 521: 	240 
    -- CP-element group 521: 	247 
    -- CP-element group 521: 	219 
    -- CP-element group 521: 	254 
    -- CP-element group 521: 	226 
    -- CP-element group 521: 	233 
    -- CP-element group 521: 	257 
    -- CP-element group 521: 	212 
    -- CP-element group 521:  members (56) 
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/addr_of_538_complete/$entry
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_548_update_start_
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_final_index_sum_regn_update_start
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_541_sample_start_
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_548_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_548_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_33/merge_stmt_524__exit__
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711__entry__
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/addr_of_538_complete/req
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_index_scale_1/scale_rename_ack
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_index_resize_1/index_resize_req
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_index_resize_1/$exit
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_index_resize_1/$entry
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_index_computed_1
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_index_scale_1/scale_rename_req
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_index_scaled_1
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_index_scale_1/$exit
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_index_resized_1
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_index_scale_1/$entry
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_final_index_sum_regn_Update/req
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_final_index_sum_regn_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_541_Sample/rr
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_final_index_sum_regn_Sample/req
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_index_resize_1/index_resize_ack
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/addr_of_538_update_start_
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/RPIPE_ConvTranspose_input_pipe_541_Sample/$entry
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/$entry
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/array_obj_ref_537_final_index_sum_regn_Sample/$entry
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_564_update_start_
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_564_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_564_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_585_update_start_
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_585_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_585_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_606_update_start_
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_606_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_606_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_627_update_start_
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_627_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_627_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_648_update_start_
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_648_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_648_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_669_update_start_
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_669_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_669_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_690_update_start_
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_690_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/type_cast_690_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_update_start_
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_Update/word_access_complete/$entry
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_Update/word_access_complete/word_0/$entry
      -- CP-element group 521: 	 branch_block_stmt_33/assign_stmt_539_to_assign_stmt_711/ptr_deref_698_Update/word_access_complete/word_0/cr
      -- CP-element group 521: 	 branch_block_stmt_33/merge_stmt_524_PhiAck/$exit
      -- CP-element group 521: 	 branch_block_stmt_33/merge_stmt_524_PhiAck/phi_stmt_525_ack
      -- 
    phi_stmt_525_ack_3672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 521_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_525_ack_0, ack => convTranspose_CP_39_elements(521)); -- 
    cr_1379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(521), ack => type_cast_548_inst_req_1); -- 
    req_1337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(521), ack => addr_of_538_final_reg_req_1); -- 
    req_1322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(521), ack => array_obj_ref_537_index_offset_req_1); -- 
    rr_1346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(521), ack => RPIPE_ConvTranspose_input_pipe_541_inst_req_0); -- 
    req_1317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(521), ack => array_obj_ref_537_index_offset_req_0); -- 
    cr_1421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(521), ack => type_cast_564_inst_req_1); -- 
    cr_1463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(521), ack => type_cast_585_inst_req_1); -- 
    cr_1505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(521), ack => type_cast_606_inst_req_1); -- 
    cr_1547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(521), ack => type_cast_627_inst_req_1); -- 
    cr_1589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(521), ack => type_cast_648_inst_req_1); -- 
    cr_1631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(521), ack => type_cast_669_inst_req_1); -- 
    cr_1673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(521), ack => type_cast_690_inst_req_1); -- 
    cr_1723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(521), ack => ptr_deref_698_store_0_req_1); -- 
    -- CP-element group 522:  transition  output  delay-element  bypass 
    -- CP-element group 522: predecessors 
    -- CP-element group 522: 	262 
    -- CP-element group 522: successors 
    -- CP-element group 522: 	526 
    -- CP-element group 522:  members (5) 
      -- CP-element group 522: 	 branch_block_stmt_33/bbx_xnph573_forx_xbody308_PhiReq/$exit
      -- CP-element group 522: 	 branch_block_stmt_33/bbx_xnph573_forx_xbody308_PhiReq/phi_stmt_756/$exit
      -- CP-element group 522: 	 branch_block_stmt_33/bbx_xnph573_forx_xbody308_PhiReq/phi_stmt_756/phi_stmt_756_sources/$exit
      -- CP-element group 522: 	 branch_block_stmt_33/bbx_xnph573_forx_xbody308_PhiReq/phi_stmt_756/phi_stmt_756_sources/type_cast_760_konst_delay_trans
      -- CP-element group 522: 	 branch_block_stmt_33/bbx_xnph573_forx_xbody308_PhiReq/phi_stmt_756/phi_stmt_756_req
      -- 
    phi_stmt_756_req_3695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_756_req_3695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(522), ack => phi_stmt_756_req_0); -- 
    -- Element group convTranspose_CP_39_elements(522) is a control-delay.
    cp_element_522_delay: control_delay_element  generic map(name => " 522_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(262), ack => convTranspose_CP_39_elements(522), clk => clk, reset =>reset);
    -- CP-element group 523:  transition  input  bypass 
    -- CP-element group 523: predecessors 
    -- CP-element group 523: 	327 
    -- CP-element group 523: successors 
    -- CP-element group 523: 	525 
    -- CP-element group 523:  members (2) 
      -- CP-element group 523: 	 branch_block_stmt_33/forx_xbody308_forx_xbody308_PhiReq/phi_stmt_756/phi_stmt_756_sources/type_cast_762/SplitProtocol/Sample/$exit
      -- CP-element group 523: 	 branch_block_stmt_33/forx_xbody308_forx_xbody308_PhiReq/phi_stmt_756/phi_stmt_756_sources/type_cast_762/SplitProtocol/Sample/ra
      -- 
    ra_3715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 523_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_762_inst_ack_0, ack => convTranspose_CP_39_elements(523)); -- 
    -- CP-element group 524:  transition  input  bypass 
    -- CP-element group 524: predecessors 
    -- CP-element group 524: 	327 
    -- CP-element group 524: successors 
    -- CP-element group 524: 	525 
    -- CP-element group 524:  members (2) 
      -- CP-element group 524: 	 branch_block_stmt_33/forx_xbody308_forx_xbody308_PhiReq/phi_stmt_756/phi_stmt_756_sources/type_cast_762/SplitProtocol/Update/$exit
      -- CP-element group 524: 	 branch_block_stmt_33/forx_xbody308_forx_xbody308_PhiReq/phi_stmt_756/phi_stmt_756_sources/type_cast_762/SplitProtocol/Update/ca
      -- 
    ca_3720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 524_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_762_inst_ack_1, ack => convTranspose_CP_39_elements(524)); -- 
    -- CP-element group 525:  join  transition  output  bypass 
    -- CP-element group 525: predecessors 
    -- CP-element group 525: 	523 
    -- CP-element group 525: 	524 
    -- CP-element group 525: successors 
    -- CP-element group 525: 	526 
    -- CP-element group 525:  members (6) 
      -- CP-element group 525: 	 branch_block_stmt_33/forx_xbody308_forx_xbody308_PhiReq/$exit
      -- CP-element group 525: 	 branch_block_stmt_33/forx_xbody308_forx_xbody308_PhiReq/phi_stmt_756/$exit
      -- CP-element group 525: 	 branch_block_stmt_33/forx_xbody308_forx_xbody308_PhiReq/phi_stmt_756/phi_stmt_756_sources/$exit
      -- CP-element group 525: 	 branch_block_stmt_33/forx_xbody308_forx_xbody308_PhiReq/phi_stmt_756/phi_stmt_756_sources/type_cast_762/$exit
      -- CP-element group 525: 	 branch_block_stmt_33/forx_xbody308_forx_xbody308_PhiReq/phi_stmt_756/phi_stmt_756_sources/type_cast_762/SplitProtocol/$exit
      -- CP-element group 525: 	 branch_block_stmt_33/forx_xbody308_forx_xbody308_PhiReq/phi_stmt_756/phi_stmt_756_req
      -- 
    phi_stmt_756_req_3721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_756_req_3721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(525), ack => phi_stmt_756_req_1); -- 
    convTranspose_cp_element_group_525: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_525"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(523) & convTranspose_CP_39_elements(524);
      gj_convTranspose_cp_element_group_525 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(525), clk => clk, reset => reset); --
    end block;
    -- CP-element group 526:  merge  transition  place  bypass 
    -- CP-element group 526: predecessors 
    -- CP-element group 526: 	525 
    -- CP-element group 526: 	522 
    -- CP-element group 526: successors 
    -- CP-element group 526: 	527 
    -- CP-element group 526:  members (2) 
      -- CP-element group 526: 	 branch_block_stmt_33/merge_stmt_755_PhiReqMerge
      -- CP-element group 526: 	 branch_block_stmt_33/merge_stmt_755_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(526) <= OrReduce(convTranspose_CP_39_elements(525) & convTranspose_CP_39_elements(522));
    -- CP-element group 527:  fork  transition  place  input  output  bypass 
    -- CP-element group 527: predecessors 
    -- CP-element group 527: 	526 
    -- CP-element group 527: successors 
    -- CP-element group 527: 	300 
    -- CP-element group 527: 	307 
    -- CP-element group 527: 	314 
    -- CP-element group 527: 	321 
    -- CP-element group 527: 	324 
    -- CP-element group 527: 	263 
    -- CP-element group 527: 	264 
    -- CP-element group 527: 	266 
    -- CP-element group 527: 	267 
    -- CP-element group 527: 	272 
    -- CP-element group 527: 	279 
    -- CP-element group 527: 	286 
    -- CP-element group 527: 	293 
    -- CP-element group 527:  members (56) 
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_921_update_start_
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_921_Update/cr
      -- CP-element group 527: 	 branch_block_stmt_33/merge_stmt_755__exit__
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942__entry__
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_858_update_start_
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_816_update_start_
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_816_Update/cr
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_921_Update/$entry
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_900_Update/$entry
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_900_Update/cr
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_858_Update/$entry
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_900_update_start_
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_Update/word_access_complete/word_0/cr
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_858_Update/cr
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_Update/word_access_complete/word_0/$entry
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_Update/word_access_complete/$entry
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_Update/$entry
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_837_Update/cr
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_837_Update/$entry
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_837_update_start_
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/ptr_deref_929_update_start_
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_879_Update/cr
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_816_Update/$entry
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_879_Update/$entry
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_879_update_start_
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/$entry
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/addr_of_769_update_start_
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_index_resized_1
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_index_scaled_1
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_index_computed_1
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_index_resize_1/$entry
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_index_resize_1/$exit
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_index_resize_1/index_resize_req
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_index_resize_1/index_resize_ack
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_index_scale_1/$entry
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_index_scale_1/$exit
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_index_scale_1/scale_rename_req
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_index_scale_1/scale_rename_ack
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_final_index_sum_regn_update_start
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_final_index_sum_regn_Sample/$entry
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_final_index_sum_regn_Sample/req
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_final_index_sum_regn_Update/$entry
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/array_obj_ref_768_final_index_sum_regn_Update/req
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/addr_of_769_complete/$entry
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/addr_of_769_complete/req
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_772_sample_start_
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_772_Sample/$entry
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/RPIPE_ConvTranspose_input_pipe_772_Sample/rr
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_779_update_start_
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_779_Update/$entry
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_779_Update/cr
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_795_update_start_
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_795_Update/$entry
      -- CP-element group 527: 	 branch_block_stmt_33/assign_stmt_770_to_assign_stmt_942/type_cast_795_Update/cr
      -- CP-element group 527: 	 branch_block_stmt_33/merge_stmt_755_PhiAck/$exit
      -- CP-element group 527: 	 branch_block_stmt_33/merge_stmt_755_PhiAck/phi_stmt_756_ack
      -- 
    phi_stmt_756_ack_3726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 527_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_756_ack_0, ack => convTranspose_CP_39_elements(527)); -- 
    cr_2144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(527), ack => type_cast_921_inst_req_1); -- 
    cr_1934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(527), ack => type_cast_816_inst_req_1); -- 
    cr_2102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(527), ack => type_cast_900_inst_req_1); -- 
    cr_2194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(527), ack => ptr_deref_929_store_0_req_1); -- 
    cr_2018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(527), ack => type_cast_858_inst_req_1); -- 
    cr_1976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(527), ack => type_cast_837_inst_req_1); -- 
    cr_2060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(527), ack => type_cast_879_inst_req_1); -- 
    req_1788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(527), ack => array_obj_ref_768_index_offset_req_0); -- 
    req_1793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(527), ack => array_obj_ref_768_index_offset_req_1); -- 
    req_1808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(527), ack => addr_of_769_final_reg_req_1); -- 
    rr_1817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(527), ack => RPIPE_ConvTranspose_input_pipe_772_inst_req_0); -- 
    cr_1850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(527), ack => type_cast_779_inst_req_1); -- 
    cr_1892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(527), ack => type_cast_795_inst_req_1); -- 
    -- CP-element group 528:  merge  fork  transition  place  output  bypass 
    -- CP-element group 528: predecessors 
    -- CP-element group 528: 	326 
    -- CP-element group 528: 	193 
    -- CP-element group 528: successors 
    -- CP-element group 528: 	328 
    -- CP-element group 528: 	329 
    -- CP-element group 528: 	330 
    -- CP-element group 528: 	331 
    -- CP-element group 528: 	332 
    -- CP-element group 528: 	333 
    -- CP-element group 528:  members (25) 
      -- CP-element group 528: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_962_Update/$entry
      -- CP-element group 528: 	 branch_block_stmt_33/merge_stmt_951__exit__
      -- CP-element group 528: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979__entry__
      -- CP-element group 528: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_958_Sample/rr
      -- CP-element group 528: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_958_Update/cr
      -- CP-element group 528: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_958_Update/$entry
      -- CP-element group 528: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_954_Update/$entry
      -- CP-element group 528: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_954_Update/cr
      -- CP-element group 528: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_962_Update/cr
      -- CP-element group 528: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_958_sample_start_
      -- CP-element group 528: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_954_Sample/rr
      -- CP-element group 528: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_954_Sample/$entry
      -- CP-element group 528: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_954_update_start_
      -- CP-element group 528: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_954_sample_start_
      -- CP-element group 528: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_958_Sample/$entry
      -- CP-element group 528: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_962_Sample/rr
      -- CP-element group 528: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/$entry
      -- CP-element group 528: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_962_Sample/$entry
      -- CP-element group 528: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_962_update_start_
      -- CP-element group 528: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_958_update_start_
      -- CP-element group 528: 	 branch_block_stmt_33/assign_stmt_955_to_assign_stmt_979/type_cast_962_sample_start_
      -- CP-element group 528: 	 branch_block_stmt_33/merge_stmt_951_PhiReqMerge
      -- CP-element group 528: 	 branch_block_stmt_33/merge_stmt_951_PhiAck/$entry
      -- CP-element group 528: 	 branch_block_stmt_33/merge_stmt_951_PhiAck/$exit
      -- CP-element group 528: 	 branch_block_stmt_33/merge_stmt_951_PhiAck/dummy
      -- 
    rr_2239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => type_cast_958_inst_req_0); -- 
    cr_2244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => type_cast_958_inst_req_1); -- 
    cr_2230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => type_cast_954_inst_req_1); -- 
    cr_2258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => type_cast_962_inst_req_1); -- 
    rr_2225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => type_cast_954_inst_req_0); -- 
    rr_2253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => type_cast_962_inst_req_0); -- 
    convTranspose_CP_39_elements(528) <= OrReduce(convTranspose_CP_39_elements(326) & convTranspose_CP_39_elements(193));
    -- CP-element group 529:  transition  output  delay-element  bypass 
    -- CP-element group 529: predecessors 
    -- CP-element group 529: 	338 
    -- CP-element group 529: successors 
    -- CP-element group 529: 	533 
    -- CP-element group 529:  members (5) 
      -- CP-element group 529: 	 branch_block_stmt_33/bbx_xnph569_forx_xbody410_PhiReq/$exit
      -- CP-element group 529: 	 branch_block_stmt_33/bbx_xnph569_forx_xbody410_PhiReq/phi_stmt_1024/$exit
      -- CP-element group 529: 	 branch_block_stmt_33/bbx_xnph569_forx_xbody410_PhiReq/phi_stmt_1024/phi_stmt_1024_sources/$exit
      -- CP-element group 529: 	 branch_block_stmt_33/bbx_xnph569_forx_xbody410_PhiReq/phi_stmt_1024/phi_stmt_1024_sources/type_cast_1028_konst_delay_trans
      -- CP-element group 529: 	 branch_block_stmt_33/bbx_xnph569_forx_xbody410_PhiReq/phi_stmt_1024/phi_stmt_1024_req
      -- 
    phi_stmt_1024_req_3772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1024_req_3772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(529), ack => phi_stmt_1024_req_0); -- 
    -- Element group convTranspose_CP_39_elements(529) is a control-delay.
    cp_element_529_delay: control_delay_element  generic map(name => " 529_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(338), ack => convTranspose_CP_39_elements(529), clk => clk, reset =>reset);
    -- CP-element group 530:  transition  input  bypass 
    -- CP-element group 530: predecessors 
    -- CP-element group 530: 	347 
    -- CP-element group 530: successors 
    -- CP-element group 530: 	532 
    -- CP-element group 530:  members (2) 
      -- CP-element group 530: 	 branch_block_stmt_33/forx_xbody410_forx_xbody410_PhiReq/phi_stmt_1024/phi_stmt_1024_sources/type_cast_1030/SplitProtocol/Sample/$exit
      -- CP-element group 530: 	 branch_block_stmt_33/forx_xbody410_forx_xbody410_PhiReq/phi_stmt_1024/phi_stmt_1024_sources/type_cast_1030/SplitProtocol/Sample/ra
      -- 
    ra_3792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 530_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1030_inst_ack_0, ack => convTranspose_CP_39_elements(530)); -- 
    -- CP-element group 531:  transition  input  bypass 
    -- CP-element group 531: predecessors 
    -- CP-element group 531: 	347 
    -- CP-element group 531: successors 
    -- CP-element group 531: 	532 
    -- CP-element group 531:  members (2) 
      -- CP-element group 531: 	 branch_block_stmt_33/forx_xbody410_forx_xbody410_PhiReq/phi_stmt_1024/phi_stmt_1024_sources/type_cast_1030/SplitProtocol/Update/$exit
      -- CP-element group 531: 	 branch_block_stmt_33/forx_xbody410_forx_xbody410_PhiReq/phi_stmt_1024/phi_stmt_1024_sources/type_cast_1030/SplitProtocol/Update/ca
      -- 
    ca_3797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 531_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1030_inst_ack_1, ack => convTranspose_CP_39_elements(531)); -- 
    -- CP-element group 532:  join  transition  output  bypass 
    -- CP-element group 532: predecessors 
    -- CP-element group 532: 	530 
    -- CP-element group 532: 	531 
    -- CP-element group 532: successors 
    -- CP-element group 532: 	533 
    -- CP-element group 532:  members (6) 
      -- CP-element group 532: 	 branch_block_stmt_33/forx_xbody410_forx_xbody410_PhiReq/$exit
      -- CP-element group 532: 	 branch_block_stmt_33/forx_xbody410_forx_xbody410_PhiReq/phi_stmt_1024/$exit
      -- CP-element group 532: 	 branch_block_stmt_33/forx_xbody410_forx_xbody410_PhiReq/phi_stmt_1024/phi_stmt_1024_sources/$exit
      -- CP-element group 532: 	 branch_block_stmt_33/forx_xbody410_forx_xbody410_PhiReq/phi_stmt_1024/phi_stmt_1024_sources/type_cast_1030/$exit
      -- CP-element group 532: 	 branch_block_stmt_33/forx_xbody410_forx_xbody410_PhiReq/phi_stmt_1024/phi_stmt_1024_sources/type_cast_1030/SplitProtocol/$exit
      -- CP-element group 532: 	 branch_block_stmt_33/forx_xbody410_forx_xbody410_PhiReq/phi_stmt_1024/phi_stmt_1024_req
      -- 
    phi_stmt_1024_req_3798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1024_req_3798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(532), ack => phi_stmt_1024_req_1); -- 
    convTranspose_cp_element_group_532: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_532"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(530) & convTranspose_CP_39_elements(531);
      gj_convTranspose_cp_element_group_532 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(532), clk => clk, reset => reset); --
    end block;
    -- CP-element group 533:  merge  transition  place  bypass 
    -- CP-element group 533: predecessors 
    -- CP-element group 533: 	529 
    -- CP-element group 533: 	532 
    -- CP-element group 533: successors 
    -- CP-element group 533: 	534 
    -- CP-element group 533:  members (2) 
      -- CP-element group 533: 	 branch_block_stmt_33/merge_stmt_1023_PhiReqMerge
      -- CP-element group 533: 	 branch_block_stmt_33/merge_stmt_1023_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(533) <= OrReduce(convTranspose_CP_39_elements(529) & convTranspose_CP_39_elements(532));
    -- CP-element group 534:  fork  transition  place  input  output  bypass 
    -- CP-element group 534: predecessors 
    -- CP-element group 534: 	533 
    -- CP-element group 534: successors 
    -- CP-element group 534: 	339 
    -- CP-element group 534: 	340 
    -- CP-element group 534: 	342 
    -- CP-element group 534: 	344 
    -- CP-element group 534:  members (29) 
      -- CP-element group 534: 	 branch_block_stmt_33/merge_stmt_1023__exit__
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054__entry__
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_final_index_sum_regn_Update/req
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_final_index_sum_regn_Update/$entry
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_final_index_sum_regn_Sample/req
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_final_index_sum_regn_Sample/$entry
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_final_index_sum_regn_update_start
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_index_scale_1/scale_rename_ack
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_index_scale_1/scale_rename_req
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_index_scale_1/$exit
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_index_scale_1/$entry
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_index_resize_1/index_resize_ack
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_index_resize_1/index_resize_req
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/addr_of_1037_complete/req
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_index_resize_1/$exit
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_index_resize_1/$entry
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/addr_of_1037_complete/$entry
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_index_computed_1
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_index_scaled_1
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/array_obj_ref_1036_index_resized_1
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_update_start_
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/addr_of_1037_update_start_
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/$entry
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_Update/$entry
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_Update/word_access_complete/$entry
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_Update/word_access_complete/word_0/$entry
      -- CP-element group 534: 	 branch_block_stmt_33/assign_stmt_1038_to_assign_stmt_1054/ptr_deref_1040_Update/word_access_complete/word_0/cr
      -- CP-element group 534: 	 branch_block_stmt_33/merge_stmt_1023_PhiAck/$exit
      -- CP-element group 534: 	 branch_block_stmt_33/merge_stmt_1023_PhiAck/phi_stmt_1024_ack
      -- 
    phi_stmt_1024_ack_3803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 534_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1024_ack_0, ack => convTranspose_CP_39_elements(534)); -- 
    req_2328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(534), ack => array_obj_ref_1036_index_offset_req_1); -- 
    req_2323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(534), ack => array_obj_ref_1036_index_offset_req_0); -- 
    req_2343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(534), ack => addr_of_1037_final_reg_req_1); -- 
    cr_2393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(534), ack => ptr_deref_1040_store_0_req_1); -- 
    -- CP-element group 535:  merge  fork  transition  place  output  bypass 
    -- CP-element group 535: predecessors 
    -- CP-element group 535: 	336 
    -- CP-element group 535: 	346 
    -- CP-element group 535: successors 
    -- CP-element group 535: 	348 
    -- CP-element group 535: 	349 
    -- CP-element group 535: 	351 
    -- CP-element group 535: 	352 
    -- CP-element group 535: 	376 
    -- CP-element group 535: 	424 
    -- CP-element group 535: 	448 
    -- CP-element group 535: 	450 
    -- CP-element group 535: 	452 
    -- CP-element group 535: 	454 
    -- CP-element group 535: 	400 
    -- CP-element group 535:  members (40) 
      -- CP-element group 535: 	 branch_block_stmt_33/merge_stmt_1063__exit__
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228__entry__
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block3_done_1227_Sample/rr
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block3_done_1227_Sample/$entry
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block3_done_1227_sample_start_
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block2_done_1224_Sample/rr
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block2_done_1224_Sample/$entry
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/$entry
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/call_stmt_1066_sample_start_
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/call_stmt_1066_update_start_
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/call_stmt_1066_Sample/$entry
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/call_stmt_1066_Sample/crr
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/call_stmt_1066_Update/$entry
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/call_stmt_1066_Update/ccr
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/type_cast_1071_update_start_
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/type_cast_1071_Update/$entry
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/type_cast_1071_Update/cr
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1073_sample_start_
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block2_done_1224_sample_start_
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1073_Sample/$entry
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block0_start_1073_Sample/req
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block1_done_1221_Sample/rr
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block1_done_1221_Sample/$entry
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block1_done_1221_sample_start_
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block0_done_1218_Sample/rr
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block0_done_1218_Sample/$entry
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/RPIPE_Block0_done_1218_sample_start_
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1109_sample_start_
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1109_Sample/$entry
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block1_start_1109_Sample/req
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1145_sample_start_
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1145_Sample/$entry
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block2_start_1145_Sample/req
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1181_sample_start_
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1181_Sample/$entry
      -- CP-element group 535: 	 branch_block_stmt_33/call_stmt_1066_to_assign_stmt_1228/WPIPE_Block3_start_1181_Sample/req
      -- CP-element group 535: 	 branch_block_stmt_33/merge_stmt_1063_PhiReqMerge
      -- CP-element group 535: 	 branch_block_stmt_33/merge_stmt_1063_PhiAck/$entry
      -- CP-element group 535: 	 branch_block_stmt_33/merge_stmt_1063_PhiAck/$exit
      -- CP-element group 535: 	 branch_block_stmt_33/merge_stmt_1063_PhiAck/dummy
      -- 
    rr_3166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(535), ack => RPIPE_Block3_done_1227_inst_req_0); -- 
    rr_3152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(535), ack => RPIPE_Block2_done_1224_inst_req_0); -- 
    crr_2424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(535), ack => call_stmt_1066_call_req_0); -- 
    ccr_2429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(535), ack => call_stmt_1066_call_req_1); -- 
    cr_2443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(535), ack => type_cast_1071_inst_req_1); -- 
    req_2452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(535), ack => WPIPE_Block0_start_1073_inst_req_0); -- 
    rr_3138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(535), ack => RPIPE_Block1_done_1221_inst_req_0); -- 
    rr_3124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(535), ack => RPIPE_Block0_done_1218_inst_req_0); -- 
    req_2620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(535), ack => WPIPE_Block1_start_1109_inst_req_0); -- 
    req_2788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(535), ack => WPIPE_Block2_start_1145_inst_req_0); -- 
    req_2956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(535), ack => WPIPE_Block3_start_1181_inst_req_0); -- 
    convTranspose_CP_39_elements(535) <= OrReduce(convTranspose_CP_39_elements(336) & convTranspose_CP_39_elements(346));
    -- CP-element group 536:  transition  output  delay-element  bypass 
    -- CP-element group 536: predecessors 
    -- CP-element group 536: 	466 
    -- CP-element group 536: successors 
    -- CP-element group 536: 	540 
    -- CP-element group 536:  members (5) 
      -- CP-element group 536: 	 branch_block_stmt_33/bbx_xnph_forx_xbody490_PhiReq/$exit
      -- CP-element group 536: 	 branch_block_stmt_33/bbx_xnph_forx_xbody490_PhiReq/phi_stmt_1290/$exit
      -- CP-element group 536: 	 branch_block_stmt_33/bbx_xnph_forx_xbody490_PhiReq/phi_stmt_1290/phi_stmt_1290_sources/$exit
      -- CP-element group 536: 	 branch_block_stmt_33/bbx_xnph_forx_xbody490_PhiReq/phi_stmt_1290/phi_stmt_1290_sources/type_cast_1296_konst_delay_trans
      -- CP-element group 536: 	 branch_block_stmt_33/bbx_xnph_forx_xbody490_PhiReq/phi_stmt_1290/phi_stmt_1290_req
      -- 
    phi_stmt_1290_req_3849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1290_req_3849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(536), ack => phi_stmt_1290_req_1); -- 
    -- Element group convTranspose_CP_39_elements(536) is a control-delay.
    cp_element_536_delay: control_delay_element  generic map(name => " 536_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(466), ack => convTranspose_CP_39_elements(536), clk => clk, reset =>reset);
    -- CP-element group 537:  transition  input  bypass 
    -- CP-element group 537: predecessors 
    -- CP-element group 537: 	514 
    -- CP-element group 537: successors 
    -- CP-element group 537: 	539 
    -- CP-element group 537:  members (2) 
      -- CP-element group 537: 	 branch_block_stmt_33/forx_xbody490_forx_xbody490_PhiReq/phi_stmt_1290/phi_stmt_1290_sources/type_cast_1293/SplitProtocol/Sample/$exit
      -- CP-element group 537: 	 branch_block_stmt_33/forx_xbody490_forx_xbody490_PhiReq/phi_stmt_1290/phi_stmt_1290_sources/type_cast_1293/SplitProtocol/Sample/ra
      -- 
    ra_3869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 537_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1293_inst_ack_0, ack => convTranspose_CP_39_elements(537)); -- 
    -- CP-element group 538:  transition  input  bypass 
    -- CP-element group 538: predecessors 
    -- CP-element group 538: 	514 
    -- CP-element group 538: successors 
    -- CP-element group 538: 	539 
    -- CP-element group 538:  members (2) 
      -- CP-element group 538: 	 branch_block_stmt_33/forx_xbody490_forx_xbody490_PhiReq/phi_stmt_1290/phi_stmt_1290_sources/type_cast_1293/SplitProtocol/Update/$exit
      -- CP-element group 538: 	 branch_block_stmt_33/forx_xbody490_forx_xbody490_PhiReq/phi_stmt_1290/phi_stmt_1290_sources/type_cast_1293/SplitProtocol/Update/ca
      -- 
    ca_3874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 538_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1293_inst_ack_1, ack => convTranspose_CP_39_elements(538)); -- 
    -- CP-element group 539:  join  transition  output  bypass 
    -- CP-element group 539: predecessors 
    -- CP-element group 539: 	538 
    -- CP-element group 539: 	537 
    -- CP-element group 539: successors 
    -- CP-element group 539: 	540 
    -- CP-element group 539:  members (6) 
      -- CP-element group 539: 	 branch_block_stmt_33/forx_xbody490_forx_xbody490_PhiReq/$exit
      -- CP-element group 539: 	 branch_block_stmt_33/forx_xbody490_forx_xbody490_PhiReq/phi_stmt_1290/$exit
      -- CP-element group 539: 	 branch_block_stmt_33/forx_xbody490_forx_xbody490_PhiReq/phi_stmt_1290/phi_stmt_1290_sources/$exit
      -- CP-element group 539: 	 branch_block_stmt_33/forx_xbody490_forx_xbody490_PhiReq/phi_stmt_1290/phi_stmt_1290_sources/type_cast_1293/$exit
      -- CP-element group 539: 	 branch_block_stmt_33/forx_xbody490_forx_xbody490_PhiReq/phi_stmt_1290/phi_stmt_1290_sources/type_cast_1293/SplitProtocol/$exit
      -- CP-element group 539: 	 branch_block_stmt_33/forx_xbody490_forx_xbody490_PhiReq/phi_stmt_1290/phi_stmt_1290_req
      -- 
    phi_stmt_1290_req_3875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1290_req_3875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(539), ack => phi_stmt_1290_req_0); -- 
    convTranspose_cp_element_group_539: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_539"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(538) & convTranspose_CP_39_elements(537);
      gj_convTranspose_cp_element_group_539 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(539), clk => clk, reset => reset); --
    end block;
    -- CP-element group 540:  merge  transition  place  bypass 
    -- CP-element group 540: predecessors 
    -- CP-element group 540: 	539 
    -- CP-element group 540: 	536 
    -- CP-element group 540: successors 
    -- CP-element group 540: 	541 
    -- CP-element group 540:  members (2) 
      -- CP-element group 540: 	 branch_block_stmt_33/merge_stmt_1289_PhiReqMerge
      -- CP-element group 540: 	 branch_block_stmt_33/merge_stmt_1289_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(540) <= OrReduce(convTranspose_CP_39_elements(539) & convTranspose_CP_39_elements(536));
    -- CP-element group 541:  fork  transition  place  input  output  bypass 
    -- CP-element group 541: predecessors 
    -- CP-element group 541: 	540 
    -- CP-element group 541: successors 
    -- CP-element group 541: 	474 
    -- CP-element group 541: 	476 
    -- CP-element group 541: 	478 
    -- CP-element group 541: 	470 
    -- CP-element group 541: 	472 
    -- CP-element group 541: 	480 
    -- CP-element group 541: 	482 
    -- CP-element group 541: 	484 
    -- CP-element group 541: 	467 
    -- CP-element group 541: 	468 
    -- CP-element group 541: 	486 
    -- CP-element group 541: 	488 
    -- CP-element group 541:  members (53) 
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/addr_of_1303_complete/$entry
      -- CP-element group 541: 	 branch_block_stmt_33/merge_stmt_1289__exit__
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417__entry__
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/addr_of_1303_update_start_
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/$entry
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_final_index_sum_regn_Sample/req
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_index_resized_1
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/addr_of_1303_complete/req
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_index_scaled_1
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_index_computed_1
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_final_index_sum_regn_Update/$entry
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_final_index_sum_regn_Update/req
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_index_resize_1/$entry
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_index_resize_1/$exit
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_index_resize_1/index_resize_req
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_index_resize_1/index_resize_ack
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_index_scale_1/$entry
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_index_scale_1/$exit
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_index_scale_1/scale_rename_req
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_final_index_sum_regn_Sample/$entry
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_final_index_sum_regn_update_start
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_update_start_
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/array_obj_ref_1302_index_scale_1/scale_rename_ack
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_Update/word_access_complete/word_0/cr
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_Update/word_access_complete/word_0/$entry
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_Update/word_access_complete/$entry
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/ptr_deref_1307_Update/$entry
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1311_update_start_
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1311_Update/$entry
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1311_Update/cr
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1321_update_start_
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1321_Update/$entry
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1321_Update/cr
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1331_update_start_
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1331_Update/$entry
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1331_Update/cr
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1341_update_start_
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1341_Update/$entry
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1341_Update/cr
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1351_update_start_
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1351_Update/$entry
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1351_Update/cr
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1361_update_start_
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1361_Update/$entry
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1361_Update/cr
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1371_update_start_
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1371_Update/$entry
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1371_Update/cr
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1381_update_start_
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1381_Update/$entry
      -- CP-element group 541: 	 branch_block_stmt_33/assign_stmt_1304_to_assign_stmt_1417/type_cast_1381_Update/cr
      -- CP-element group 541: 	 branch_block_stmt_33/merge_stmt_1289_PhiAck/$exit
      -- CP-element group 541: 	 branch_block_stmt_33/merge_stmt_1289_PhiAck/phi_stmt_1290_ack
      -- 
    phi_stmt_1290_ack_3880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 541_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1290_ack_0, ack => convTranspose_CP_39_elements(541)); -- 
    req_3281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(541), ack => array_obj_ref_1302_index_offset_req_0); -- 
    req_3301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(541), ack => addr_of_1303_final_reg_req_1); -- 
    req_3286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(541), ack => array_obj_ref_1302_index_offset_req_1); -- 
    cr_3346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(541), ack => ptr_deref_1307_load_0_req_1); -- 
    cr_3365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(541), ack => type_cast_1311_inst_req_1); -- 
    cr_3379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(541), ack => type_cast_1321_inst_req_1); -- 
    cr_3393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(541), ack => type_cast_1331_inst_req_1); -- 
    cr_3407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(541), ack => type_cast_1341_inst_req_1); -- 
    cr_3421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(541), ack => type_cast_1351_inst_req_1); -- 
    cr_3435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(541), ack => type_cast_1361_inst_req_1); -- 
    cr_3449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(541), ack => type_cast_1371_inst_req_1); -- 
    cr_3463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(541), ack => type_cast_1381_inst_req_1); -- 
    -- CP-element group 542:  merge  transition  place  bypass 
    -- CP-element group 542: predecessors 
    -- CP-element group 542: 	513 
    -- CP-element group 542: 	464 
    -- CP-element group 542: successors 
    -- CP-element group 542:  members (16) 
      -- CP-element group 542: 	 $exit
      -- CP-element group 542: 	 branch_block_stmt_33/$exit
      -- CP-element group 542: 	 branch_block_stmt_33/branch_block_stmt_33__exit__
      -- CP-element group 542: 	 branch_block_stmt_33/merge_stmt_1426__exit__
      -- CP-element group 542: 	 branch_block_stmt_33/return__
      -- CP-element group 542: 	 branch_block_stmt_33/merge_stmt_1428__exit__
      -- CP-element group 542: 	 branch_block_stmt_33/merge_stmt_1426_PhiReqMerge
      -- CP-element group 542: 	 branch_block_stmt_33/merge_stmt_1426_PhiAck/$entry
      -- CP-element group 542: 	 branch_block_stmt_33/merge_stmt_1426_PhiAck/$exit
      -- CP-element group 542: 	 branch_block_stmt_33/merge_stmt_1426_PhiAck/dummy
      -- CP-element group 542: 	 branch_block_stmt_33/return___PhiReq/$entry
      -- CP-element group 542: 	 branch_block_stmt_33/return___PhiReq/$exit
      -- CP-element group 542: 	 branch_block_stmt_33/merge_stmt_1428_PhiReqMerge
      -- CP-element group 542: 	 branch_block_stmt_33/merge_stmt_1428_PhiAck/$entry
      -- CP-element group 542: 	 branch_block_stmt_33/merge_stmt_1428_PhiAck/$exit
      -- CP-element group 542: 	 branch_block_stmt_33/merge_stmt_1428_PhiAck/dummy
      -- 
    convTranspose_CP_39_elements(542) <= OrReduce(convTranspose_CP_39_elements(513) & convTranspose_CP_39_elements(464));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar587_1035_resized : std_logic_vector(13 downto 0);
    signal R_indvar587_1035_scaled : std_logic_vector(13 downto 0);
    signal R_indvar601_767_resized : std_logic_vector(10 downto 0);
    signal R_indvar601_767_scaled : std_logic_vector(10 downto 0);
    signal R_indvar617_536_resized : std_logic_vector(13 downto 0);
    signal R_indvar617_536_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1301_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1301_scaled : std_logic_vector(13 downto 0);
    signal add111_250 : std_logic_vector(15 downto 0);
    signal add148_334 : std_logic_vector(15 downto 0);
    signal add165_365 : std_logic_vector(15 downto 0);
    signal add182_396 : std_logic_vector(15 downto 0);
    signal add199_427 : std_logic_vector(15 downto 0);
    signal add216_458 : std_logic_vector(15 downto 0);
    signal add238_570 : std_logic_vector(63 downto 0);
    signal add248_591 : std_logic_vector(63 downto 0);
    signal add258_612 : std_logic_vector(63 downto 0);
    signal add268_633 : std_logic_vector(63 downto 0);
    signal add26_95 : std_logic_vector(15 downto 0);
    signal add278_654 : std_logic_vector(63 downto 0);
    signal add288_675 : std_logic_vector(63 downto 0);
    signal add298_696 : std_logic_vector(63 downto 0);
    signal add326_801 : std_logic_vector(63 downto 0);
    signal add336_822 : std_logic_vector(63 downto 0);
    signal add346_843 : std_logic_vector(63 downto 0);
    signal add356_864 : std_logic_vector(63 downto 0);
    signal add366_885 : std_logic_vector(63 downto 0);
    signal add376_906 : std_logic_vector(63 downto 0);
    signal add386_927 : std_logic_vector(63 downto 0);
    signal add43_126 : std_logic_vector(15 downto 0);
    signal add60_157 : std_logic_vector(15 downto 0);
    signal add77_188 : std_logic_vector(15 downto 0);
    signal add94_219 : std_logic_vector(15 downto 0);
    signal add_64 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1036_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1036_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1036_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1036_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1036_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1036_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1302_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1302_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1302_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1302_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1302_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1302_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_537_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_537_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_537_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_537_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_537_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_537_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_768_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_768_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_768_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_768_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_768_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_768_root_address : std_logic_vector(10 downto 0);
    signal arrayidx390_770 : std_logic_vector(31 downto 0);
    signal arrayidx413_1038 : std_logic_vector(31 downto 0);
    signal arrayidx495_1304 : std_logic_vector(31 downto 0);
    signal arrayidx_539 : std_logic_vector(31 downto 0);
    signal call107_238 : std_logic_vector(7 downto 0);
    signal call135_306 : std_logic_vector(7 downto 0);
    signal call13_67 : std_logic_vector(7 downto 0);
    signal call144_322 : std_logic_vector(7 downto 0);
    signal call152_337 : std_logic_vector(7 downto 0);
    signal call161_353 : std_logic_vector(7 downto 0);
    signal call169_368 : std_logic_vector(7 downto 0);
    signal call178_384 : std_logic_vector(7 downto 0);
    signal call186_399 : std_logic_vector(7 downto 0);
    signal call195_415 : std_logic_vector(7 downto 0);
    signal call203_430 : std_logic_vector(7 downto 0);
    signal call212_446 : std_logic_vector(7 downto 0);
    signal call225_542 : std_logic_vector(7 downto 0);
    signal call22_83 : std_logic_vector(7 downto 0);
    signal call233_558 : std_logic_vector(7 downto 0);
    signal call243_579 : std_logic_vector(7 downto 0);
    signal call253_600 : std_logic_vector(7 downto 0);
    signal call263_621 : std_logic_vector(7 downto 0);
    signal call273_642 : std_logic_vector(7 downto 0);
    signal call283_663 : std_logic_vector(7 downto 0);
    signal call293_684 : std_logic_vector(7 downto 0);
    signal call30_98 : std_logic_vector(7 downto 0);
    signal call313_773 : std_logic_vector(7 downto 0);
    signal call321_789 : std_logic_vector(7 downto 0);
    signal call331_810 : std_logic_vector(7 downto 0);
    signal call341_831 : std_logic_vector(7 downto 0);
    signal call351_852 : std_logic_vector(7 downto 0);
    signal call361_873 : std_logic_vector(7 downto 0);
    signal call371_894 : std_logic_vector(7 downto 0);
    signal call381_915 : std_logic_vector(7 downto 0);
    signal call39_114 : std_logic_vector(7 downto 0);
    signal call419_1066 : std_logic_vector(63 downto 0);
    signal call470_1219 : std_logic_vector(15 downto 0);
    signal call472_1222 : std_logic_vector(15 downto 0);
    signal call474_1225 : std_logic_vector(15 downto 0);
    signal call476_1228 : std_logic_vector(15 downto 0);
    signal call478_1231 : std_logic_vector(63 downto 0);
    signal call47_129 : std_logic_vector(7 downto 0);
    signal call56_145 : std_logic_vector(7 downto 0);
    signal call64_160 : std_logic_vector(7 downto 0);
    signal call6_52 : std_logic_vector(7 downto 0);
    signal call73_176 : std_logic_vector(7 downto 0);
    signal call81_191 : std_logic_vector(7 downto 0);
    signal call90_207 : std_logic_vector(7 downto 0);
    signal call98_222 : std_logic_vector(7 downto 0);
    signal call_36 : std_logic_vector(7 downto 0);
    signal cmp306571_480 : std_logic_vector(0 downto 0);
    signal cmp408567_979 : std_logic_vector(0 downto 0);
    signal cmp575_465 : std_logic_vector(0 downto 0);
    signal conv103_229 : std_logic_vector(15 downto 0);
    signal conv110_245 : std_logic_vector(15 downto 0);
    signal conv115_254 : std_logic_vector(31 downto 0);
    signal conv117_258 : std_logic_vector(31 downto 0);
    signal conv119_262 : std_logic_vector(31 downto 0);
    signal conv123_276 : std_logic_vector(31 downto 0);
    signal conv125_280 : std_logic_vector(31 downto 0);
    signal conv128_284 : std_logic_vector(31 downto 0);
    signal conv131_288 : std_logic_vector(31 downto 0);
    signal conv140_313 : std_logic_vector(15 downto 0);
    signal conv147_329 : std_logic_vector(15 downto 0);
    signal conv157_344 : std_logic_vector(15 downto 0);
    signal conv164_360 : std_logic_vector(15 downto 0);
    signal conv174_375 : std_logic_vector(15 downto 0);
    signal conv181_391 : std_logic_vector(15 downto 0);
    signal conv18_74 : std_logic_vector(15 downto 0);
    signal conv191_406 : std_logic_vector(15 downto 0);
    signal conv198_422 : std_logic_vector(15 downto 0);
    signal conv208_437 : std_logic_vector(15 downto 0);
    signal conv215_453 : std_logic_vector(15 downto 0);
    signal conv228_549 : std_logic_vector(63 downto 0);
    signal conv237_565 : std_logic_vector(63 downto 0);
    signal conv247_586 : std_logic_vector(63 downto 0);
    signal conv257_607 : std_logic_vector(63 downto 0);
    signal conv25_90 : std_logic_vector(15 downto 0);
    signal conv267_628 : std_logic_vector(63 downto 0);
    signal conv277_649 : std_logic_vector(63 downto 0);
    signal conv287_670 : std_logic_vector(63 downto 0);
    signal conv297_691 : std_logic_vector(63 downto 0);
    signal conv316_780 : std_logic_vector(63 downto 0);
    signal conv325_796 : std_logic_vector(63 downto 0);
    signal conv335_817 : std_logic_vector(63 downto 0);
    signal conv345_838 : std_logic_vector(63 downto 0);
    signal conv355_859 : std_logic_vector(63 downto 0);
    signal conv35_105 : std_logic_vector(15 downto 0);
    signal conv365_880 : std_logic_vector(63 downto 0);
    signal conv375_901 : std_logic_vector(63 downto 0);
    signal conv385_922 : std_logic_vector(63 downto 0);
    signal conv397_955 : std_logic_vector(31 downto 0);
    signal conv399_959 : std_logic_vector(31 downto 0);
    signal conv3_43 : std_logic_vector(15 downto 0);
    signal conv402_963 : std_logic_vector(31 downto 0);
    signal conv420_1072 : std_logic_vector(63 downto 0);
    signal conv42_121 : std_logic_vector(15 downto 0);
    signal conv479_1236 : std_logic_vector(63 downto 0);
    signal conv499_1312 : std_logic_vector(7 downto 0);
    signal conv505_1322 : std_logic_vector(7 downto 0);
    signal conv511_1332 : std_logic_vector(7 downto 0);
    signal conv517_1342 : std_logic_vector(7 downto 0);
    signal conv523_1352 : std_logic_vector(7 downto 0);
    signal conv529_1362 : std_logic_vector(7 downto 0);
    signal conv52_136 : std_logic_vector(15 downto 0);
    signal conv535_1372 : std_logic_vector(7 downto 0);
    signal conv541_1382 : std_logic_vector(7 downto 0);
    signal conv59_152 : std_logic_vector(15 downto 0);
    signal conv69_167 : std_logic_vector(15 downto 0);
    signal conv76_183 : std_logic_vector(15 downto 0);
    signal conv86_198 : std_logic_vector(15 downto 0);
    signal conv93_214 : std_logic_vector(15 downto 0);
    signal conv9_59 : std_logic_vector(15 downto 0);
    signal exitcond1_1417 : std_logic_vector(0 downto 0);
    signal exitcond2_942 : std_logic_vector(0 downto 0);
    signal exitcond3_711 : std_logic_vector(0 downto 0);
    signal exitcond_1054 : std_logic_vector(0 downto 0);
    signal iNsTr_102_740 : std_logic_vector(63 downto 0);
    signal iNsTr_132_1008 : std_logic_vector(63 downto 0);
    signal iNsTr_243_1274 : std_logic_vector(63 downto 0);
    signal iNsTr_73_509 : std_logic_vector(63 downto 0);
    signal indvar587_1024 : std_logic_vector(63 downto 0);
    signal indvar601_756 : std_logic_vector(63 downto 0);
    signal indvar617_525 : std_logic_vector(63 downto 0);
    signal indvar_1290 : std_logic_vector(63 downto 0);
    signal indvarx_xnext588_1049 : std_logic_vector(63 downto 0);
    signal indvarx_xnext602_937 : std_logic_vector(63 downto 0);
    signal indvarx_xnext618_706 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1412 : std_logic_vector(63 downto 0);
    signal mul120_272 : std_logic_vector(31 downto 0);
    signal mul126_293 : std_logic_vector(31 downto 0);
    signal mul129_298 : std_logic_vector(31 downto 0);
    signal mul132_303 : std_logic_vector(31 downto 0);
    signal mul400_968 : std_logic_vector(31 downto 0);
    signal mul403_973 : std_logic_vector(31 downto 0);
    signal mul_267 : std_logic_vector(31 downto 0);
    signal ptr_deref_1040_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1040_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1040_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1040_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1040_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1040_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1307_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1307_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1307_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1307_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1307_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_698_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_698_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_698_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_698_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_698_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_698_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_929_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_929_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_929_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_929_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_929_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_929_word_offset_0 : std_logic_vector(10 downto 0);
    signal shl104_235 : std_logic_vector(15 downto 0);
    signal shl141_319 : std_logic_vector(15 downto 0);
    signal shl158_350 : std_logic_vector(15 downto 0);
    signal shl175_381 : std_logic_vector(15 downto 0);
    signal shl192_412 : std_logic_vector(15 downto 0);
    signal shl19_80 : std_logic_vector(15 downto 0);
    signal shl209_443 : std_logic_vector(15 downto 0);
    signal shl230_555 : std_logic_vector(63 downto 0);
    signal shl240_576 : std_logic_vector(63 downto 0);
    signal shl250_597 : std_logic_vector(63 downto 0);
    signal shl260_618 : std_logic_vector(63 downto 0);
    signal shl270_639 : std_logic_vector(63 downto 0);
    signal shl280_660 : std_logic_vector(63 downto 0);
    signal shl290_681 : std_logic_vector(63 downto 0);
    signal shl318_786 : std_logic_vector(63 downto 0);
    signal shl328_807 : std_logic_vector(63 downto 0);
    signal shl338_828 : std_logic_vector(63 downto 0);
    signal shl348_849 : std_logic_vector(63 downto 0);
    signal shl358_870 : std_logic_vector(63 downto 0);
    signal shl368_891 : std_logic_vector(63 downto 0);
    signal shl36_111 : std_logic_vector(15 downto 0);
    signal shl378_912 : std_logic_vector(63 downto 0);
    signal shl53_142 : std_logic_vector(15 downto 0);
    signal shl70_173 : std_logic_vector(15 downto 0);
    signal shl87_204 : std_logic_vector(15 downto 0);
    signal shl_49 : std_logic_vector(15 downto 0);
    signal shr502_1318 : std_logic_vector(63 downto 0);
    signal shr508_1328 : std_logic_vector(63 downto 0);
    signal shr514_1338 : std_logic_vector(63 downto 0);
    signal shr520_1348 : std_logic_vector(63 downto 0);
    signal shr526_1358 : std_logic_vector(63 downto 0);
    signal shr532_1368 : std_logic_vector(63 downto 0);
    signal shr538_1378 : std_logic_vector(63 downto 0);
    signal sub_1241 : std_logic_vector(63 downto 0);
    signal tmp496_1308 : std_logic_vector(63 downto 0);
    signal tmp582_1258 : std_logic_vector(31 downto 0);
    signal tmp582x_xop_1270 : std_logic_vector(31 downto 0);
    signal tmp583_1264 : std_logic_vector(0 downto 0);
    signal tmp586_1287 : std_logic_vector(63 downto 0);
    signal tmp594_992 : std_logic_vector(31 downto 0);
    signal tmp594x_xop_1004 : std_logic_vector(31 downto 0);
    signal tmp595_998 : std_logic_vector(0 downto 0);
    signal tmp599_1021 : std_logic_vector(63 downto 0);
    signal tmp610_724 : std_logic_vector(31 downto 0);
    signal tmp610x_xop_736 : std_logic_vector(31 downto 0);
    signal tmp611_730 : std_logic_vector(0 downto 0);
    signal tmp615_753 : std_logic_vector(63 downto 0);
    signal tmp624_493 : std_logic_vector(31 downto 0);
    signal tmp624x_xop_505 : std_logic_vector(31 downto 0);
    signal tmp625_499 : std_logic_vector(0 downto 0);
    signal tmp629_522 : std_logic_vector(63 downto 0);
    signal type_cast_1002_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1012_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1019_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1028_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1030_wire : std_logic_vector(63 downto 0);
    signal type_cast_1042_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1047_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1070_wire : std_logic_vector(63 downto 0);
    signal type_cast_109_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1234_wire : std_logic_vector(63 downto 0);
    signal type_cast_1256_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1262_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1268_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1278_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1285_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1293_wire : std_logic_vector(63 downto 0);
    signal type_cast_1296_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1316_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1326_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1336_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1346_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1356_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1366_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1376_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_140_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1410_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_171_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_202_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_233_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_317_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_348_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_379_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_410_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_441_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_462_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_478_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_47_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_491_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_497_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_503_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_513_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_520_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_529_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_531_wire : std_logic_vector(63 downto 0);
    signal type_cast_553_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_574_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_595_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_616_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_637_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_658_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_679_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_704_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_722_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_728_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_734_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_744_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_751_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_760_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_762_wire : std_logic_vector(63 downto 0);
    signal type_cast_784_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_78_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_805_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_826_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_847_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_868_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_889_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_910_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_935_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_977_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_990_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_996_wire_constant : std_logic_vector(31 downto 0);
    signal xx_xop631_1014 : std_logic_vector(63 downto 0);
    signal xx_xop632_746 : std_logic_vector(63 downto 0);
    signal xx_xop633_515 : std_logic_vector(63 downto 0);
    signal xx_xop_1280 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1036_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1036_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1036_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1036_resized_base_address <= "00000000000000";
    array_obj_ref_1302_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1302_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1302_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1302_resized_base_address <= "00000000000000";
    array_obj_ref_537_constant_part_of_offset <= "00000000000000";
    array_obj_ref_537_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_537_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_537_resized_base_address <= "00000000000000";
    array_obj_ref_768_constant_part_of_offset <= "00000100010";
    array_obj_ref_768_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_768_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_768_resized_base_address <= "00000000000";
    ptr_deref_1040_word_offset_0 <= "00000000000000";
    ptr_deref_1307_word_offset_0 <= "00000000000000";
    ptr_deref_698_word_offset_0 <= "00000000000000";
    ptr_deref_929_word_offset_0 <= "00000000000";
    type_cast_1002_wire_constant <= "11111111111111111111111111111111";
    type_cast_1012_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1019_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1028_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1042_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1047_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_109_wire_constant <= "0000000000001000";
    type_cast_1256_wire_constant <= "00000000000000000000000000000010";
    type_cast_1262_wire_constant <= "00000000000000000000000000000001";
    type_cast_1268_wire_constant <= "11111111111111111111111111111111";
    type_cast_1278_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1285_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1296_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1316_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1326_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1336_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1346_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1356_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1366_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1376_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_140_wire_constant <= "0000000000001000";
    type_cast_1410_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_171_wire_constant <= "0000000000001000";
    type_cast_202_wire_constant <= "0000000000001000";
    type_cast_233_wire_constant <= "0000000000001000";
    type_cast_317_wire_constant <= "0000000000001000";
    type_cast_348_wire_constant <= "0000000000001000";
    type_cast_379_wire_constant <= "0000000000001000";
    type_cast_410_wire_constant <= "0000000000001000";
    type_cast_441_wire_constant <= "0000000000001000";
    type_cast_462_wire_constant <= "00000000000000000000000000000011";
    type_cast_478_wire_constant <= "00000000000000000000000000000011";
    type_cast_47_wire_constant <= "0000000000001000";
    type_cast_491_wire_constant <= "00000000000000000000000000000010";
    type_cast_497_wire_constant <= "00000000000000000000000000000001";
    type_cast_503_wire_constant <= "11111111111111111111111111111111";
    type_cast_513_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_520_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_529_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_553_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_574_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_595_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_616_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_637_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_658_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_679_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_704_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_722_wire_constant <= "00000000000000000000000000000010";
    type_cast_728_wire_constant <= "00000000000000000000000000000001";
    type_cast_734_wire_constant <= "11111111111111111111111111111111";
    type_cast_744_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_751_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_760_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_784_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_78_wire_constant <= "0000000000001000";
    type_cast_805_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_826_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_847_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_868_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_889_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_910_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_935_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_977_wire_constant <= "00000000000000000000000000000011";
    type_cast_990_wire_constant <= "00000000000000000000000000000010";
    type_cast_996_wire_constant <= "00000000000000000000000000000001";
    phi_stmt_1024: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1028_wire_constant & type_cast_1030_wire;
      req <= phi_stmt_1024_req_0 & phi_stmt_1024_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1024",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1024_ack_0,
          idata => idata,
          odata => indvar587_1024,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1024
    phi_stmt_1290: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1293_wire & type_cast_1296_wire_constant;
      req <= phi_stmt_1290_req_0 & phi_stmt_1290_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1290",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1290_ack_0,
          idata => idata,
          odata => indvar_1290,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1290
    phi_stmt_525: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_529_wire_constant & type_cast_531_wire;
      req <= phi_stmt_525_req_0 & phi_stmt_525_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_525",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_525_ack_0,
          idata => idata,
          odata => indvar617_525,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_525
    phi_stmt_756: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_760_wire_constant & type_cast_762_wire;
      req <= phi_stmt_756_req_0 & phi_stmt_756_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_756",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_756_ack_0,
          idata => idata,
          odata => indvar601_756,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_756
    -- flow-through select operator MUX_1020_inst
    tmp599_1021 <= xx_xop631_1014 when (tmp595_998(0) /=  '0') else type_cast_1019_wire_constant;
    -- flow-through select operator MUX_1286_inst
    tmp586_1287 <= xx_xop_1280 when (tmp583_1264(0) /=  '0') else type_cast_1285_wire_constant;
    -- flow-through select operator MUX_521_inst
    tmp629_522 <= xx_xop633_515 when (tmp625_499(0) /=  '0') else type_cast_520_wire_constant;
    -- flow-through select operator MUX_752_inst
    tmp615_753 <= xx_xop632_746 when (tmp611_730(0) /=  '0') else type_cast_751_wire_constant;
    addr_of_1037_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1037_final_reg_req_0;
      addr_of_1037_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1037_final_reg_req_1;
      addr_of_1037_final_reg_ack_1<= rack(0);
      addr_of_1037_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1037_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1036_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx413_1038,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1303_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1303_final_reg_req_0;
      addr_of_1303_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1303_final_reg_req_1;
      addr_of_1303_final_reg_ack_1<= rack(0);
      addr_of_1303_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1303_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1302_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx495_1304,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_538_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_538_final_reg_req_0;
      addr_of_538_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_538_final_reg_req_1;
      addr_of_538_final_reg_ack_1<= rack(0);
      addr_of_538_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_538_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_537_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_539,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_769_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_769_final_reg_req_0;
      addr_of_769_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_769_final_reg_req_1;
      addr_of_769_final_reg_ack_1<= rack(0);
      addr_of_769_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_769_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_768_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx390_770,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1007_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1007_inst_req_0;
      type_cast_1007_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1007_inst_req_1;
      type_cast_1007_inst_ack_1<= rack(0);
      type_cast_1007_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1007_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp594x_xop_1004,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_132_1008,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1030_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1030_inst_req_0;
      type_cast_1030_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1030_inst_req_1;
      type_cast_1030_inst_ack_1<= rack(0);
      type_cast_1030_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1030_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext588_1049,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1030_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_104_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_104_inst_req_0;
      type_cast_104_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_104_inst_req_1;
      type_cast_104_inst_ack_1<= rack(0);
      type_cast_104_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_104_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call30_98,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_105,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1071_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1071_inst_req_0;
      type_cast_1071_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1071_inst_req_1;
      type_cast_1071_inst_ack_1<= rack(0);
      type_cast_1071_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1071_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1070_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv420_1072,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_120_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_120_inst_req_0;
      type_cast_120_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_120_inst_req_1;
      type_cast_120_inst_ack_1<= rack(0);
      type_cast_120_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_120_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call39_114,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_121,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1235_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1235_inst_req_0;
      type_cast_1235_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1235_inst_req_1;
      type_cast_1235_inst_ack_1<= rack(0);
      type_cast_1235_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1235_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1234_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv479_1236,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1273_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1273_inst_req_0;
      type_cast_1273_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1273_inst_req_1;
      type_cast_1273_inst_ack_1<= rack(0);
      type_cast_1273_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1273_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp582x_xop_1270,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_243_1274,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1293_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1293_inst_req_0;
      type_cast_1293_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1293_inst_req_1;
      type_cast_1293_inst_ack_1<= rack(0);
      type_cast_1293_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1293_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1412,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1293_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1311_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1311_inst_req_0;
      type_cast_1311_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1311_inst_req_1;
      type_cast_1311_inst_ack_1<= rack(0);
      type_cast_1311_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1311_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp496_1308,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv499_1312,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1321_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1321_inst_req_0;
      type_cast_1321_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1321_inst_req_1;
      type_cast_1321_inst_ack_1<= rack(0);
      type_cast_1321_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1321_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr502_1318,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv505_1322,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1331_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1331_inst_req_0;
      type_cast_1331_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1331_inst_req_1;
      type_cast_1331_inst_ack_1<= rack(0);
      type_cast_1331_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1331_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr508_1328,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv511_1332,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1341_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1341_inst_req_0;
      type_cast_1341_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1341_inst_req_1;
      type_cast_1341_inst_ack_1<= rack(0);
      type_cast_1341_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1341_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr514_1338,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv517_1342,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1351_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1351_inst_req_0;
      type_cast_1351_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1351_inst_req_1;
      type_cast_1351_inst_ack_1<= rack(0);
      type_cast_1351_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1351_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr520_1348,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv523_1352,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_135_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_135_inst_req_0;
      type_cast_135_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_135_inst_req_1;
      type_cast_135_inst_ack_1<= rack(0);
      type_cast_135_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_135_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call47_129,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_136,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1361_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1361_inst_req_0;
      type_cast_1361_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1361_inst_req_1;
      type_cast_1361_inst_ack_1<= rack(0);
      type_cast_1361_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1361_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr526_1358,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv529_1362,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1371_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1371_inst_req_0;
      type_cast_1371_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1371_inst_req_1;
      type_cast_1371_inst_ack_1<= rack(0);
      type_cast_1371_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1371_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr532_1368,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv535_1372,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1381_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1381_inst_req_0;
      type_cast_1381_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1381_inst_req_1;
      type_cast_1381_inst_ack_1<= rack(0);
      type_cast_1381_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1381_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr538_1378,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv541_1382,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_151_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_151_inst_req_0;
      type_cast_151_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_151_inst_req_1;
      type_cast_151_inst_ack_1<= rack(0);
      type_cast_151_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_151_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call56_145,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_152,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_166_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_166_inst_req_0;
      type_cast_166_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_166_inst_req_1;
      type_cast_166_inst_ack_1<= rack(0);
      type_cast_166_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_166_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call64_160,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_167,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_182_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_182_inst_req_0;
      type_cast_182_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_182_inst_req_1;
      type_cast_182_inst_ack_1<= rack(0);
      type_cast_182_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_182_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call73_176,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv76_183,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_197_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_197_inst_req_0;
      type_cast_197_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_197_inst_req_1;
      type_cast_197_inst_ack_1<= rack(0);
      type_cast_197_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_197_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call81_191,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv86_198,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_213_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_213_inst_req_0;
      type_cast_213_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_213_inst_req_1;
      type_cast_213_inst_ack_1<= rack(0);
      type_cast_213_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_213_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call90_207,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv93_214,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_228_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_228_inst_req_0;
      type_cast_228_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_228_inst_req_1;
      type_cast_228_inst_ack_1<= rack(0);
      type_cast_228_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_228_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call98_222,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv103_229,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_244_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_244_inst_req_0;
      type_cast_244_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_244_inst_req_1;
      type_cast_244_inst_ack_1<= rack(0);
      type_cast_244_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_244_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call107_238,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv110_245,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_253_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_253_inst_req_0;
      type_cast_253_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_253_inst_req_1;
      type_cast_253_inst_ack_1<= rack(0);
      type_cast_253_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_253_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_64,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_254,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_257_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_257_inst_req_0;
      type_cast_257_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_257_inst_req_1;
      type_cast_257_inst_ack_1<= rack(0);
      type_cast_257_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_257_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add26_95,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv117_258,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_261_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_261_inst_req_0;
      type_cast_261_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_261_inst_req_1;
      type_cast_261_inst_ack_1<= rack(0);
      type_cast_261_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_261_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add43_126,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv119_262,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_275_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_275_inst_req_0;
      type_cast_275_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_275_inst_req_1;
      type_cast_275_inst_ack_1<= rack(0);
      type_cast_275_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_275_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add60_157,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv123_276,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_279_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_279_inst_req_0;
      type_cast_279_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_279_inst_req_1;
      type_cast_279_inst_ack_1<= rack(0);
      type_cast_279_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_279_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add77_188,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_280,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_283_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_283_inst_req_0;
      type_cast_283_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_283_inst_req_1;
      type_cast_283_inst_ack_1<= rack(0);
      type_cast_283_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_283_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add94_219,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv128_284,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_287_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_287_inst_req_0;
      type_cast_287_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_287_inst_req_1;
      type_cast_287_inst_ack_1<= rack(0);
      type_cast_287_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_287_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add111_250,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_288,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_312_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_312_inst_req_0;
      type_cast_312_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_312_inst_req_1;
      type_cast_312_inst_ack_1<= rack(0);
      type_cast_312_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_312_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call135_306,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv140_313,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_328_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_328_inst_req_0;
      type_cast_328_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_328_inst_req_1;
      type_cast_328_inst_ack_1<= rack(0);
      type_cast_328_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_328_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call144_322,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv147_329,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_343_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_343_inst_req_0;
      type_cast_343_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_343_inst_req_1;
      type_cast_343_inst_ack_1<= rack(0);
      type_cast_343_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_343_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call152_337,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv157_344,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_359_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_359_inst_req_0;
      type_cast_359_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_359_inst_req_1;
      type_cast_359_inst_ack_1<= rack(0);
      type_cast_359_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_359_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call161_353,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv164_360,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_374_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_374_inst_req_0;
      type_cast_374_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_374_inst_req_1;
      type_cast_374_inst_ack_1<= rack(0);
      type_cast_374_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_374_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call169_368,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv174_375,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_390_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_390_inst_req_0;
      type_cast_390_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_390_inst_req_1;
      type_cast_390_inst_ack_1<= rack(0);
      type_cast_390_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_390_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call178_384,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv181_391,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_405_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_405_inst_req_0;
      type_cast_405_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_405_inst_req_1;
      type_cast_405_inst_ack_1<= rack(0);
      type_cast_405_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_405_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call186_399,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv191_406,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_421_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_421_inst_req_0;
      type_cast_421_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_421_inst_req_1;
      type_cast_421_inst_ack_1<= rack(0);
      type_cast_421_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_421_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call195_415,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv198_422,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_42_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_42_inst_req_0;
      type_cast_42_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_42_inst_req_1;
      type_cast_42_inst_ack_1<= rack(0);
      type_cast_42_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_42_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_43,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_436_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_436_inst_req_0;
      type_cast_436_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_436_inst_req_1;
      type_cast_436_inst_ack_1<= rack(0);
      type_cast_436_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_436_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call203_430,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv208_437,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_452_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_452_inst_req_0;
      type_cast_452_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_452_inst_req_1;
      type_cast_452_inst_ack_1<= rack(0);
      type_cast_452_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_452_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call212_446,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv215_453,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_508_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_508_inst_req_0;
      type_cast_508_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_508_inst_req_1;
      type_cast_508_inst_ack_1<= rack(0);
      type_cast_508_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_508_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp624x_xop_505,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_73_509,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_531_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_531_inst_req_0;
      type_cast_531_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_531_inst_req_1;
      type_cast_531_inst_ack_1<= rack(0);
      type_cast_531_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_531_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext618_706,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_531_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_548_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_548_inst_req_0;
      type_cast_548_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_548_inst_req_1;
      type_cast_548_inst_ack_1<= rack(0);
      type_cast_548_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_548_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call225_542,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv228_549,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_564_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_564_inst_req_0;
      type_cast_564_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_564_inst_req_1;
      type_cast_564_inst_ack_1<= rack(0);
      type_cast_564_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_564_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call233_558,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv237_565,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_585_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_585_inst_req_0;
      type_cast_585_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_585_inst_req_1;
      type_cast_585_inst_ack_1<= rack(0);
      type_cast_585_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_585_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call243_579,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv247_586,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_58_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_58_inst_req_0;
      type_cast_58_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_58_inst_req_1;
      type_cast_58_inst_ack_1<= rack(0);
      type_cast_58_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_58_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_52,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9_59,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_606_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_606_inst_req_0;
      type_cast_606_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_606_inst_req_1;
      type_cast_606_inst_ack_1<= rack(0);
      type_cast_606_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_606_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call253_600,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv257_607,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_627_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_627_inst_req_0;
      type_cast_627_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_627_inst_req_1;
      type_cast_627_inst_ack_1<= rack(0);
      type_cast_627_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_627_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call263_621,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv267_628,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_648_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_648_inst_req_0;
      type_cast_648_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_648_inst_req_1;
      type_cast_648_inst_ack_1<= rack(0);
      type_cast_648_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_648_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call273_642,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv277_649,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_669_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_669_inst_req_0;
      type_cast_669_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_669_inst_req_1;
      type_cast_669_inst_ack_1<= rack(0);
      type_cast_669_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_669_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call283_663,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv287_670,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_690_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_690_inst_req_0;
      type_cast_690_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_690_inst_req_1;
      type_cast_690_inst_ack_1<= rack(0);
      type_cast_690_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_690_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call293_684,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv297_691,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_739_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_739_inst_req_0;
      type_cast_739_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_739_inst_req_1;
      type_cast_739_inst_ack_1<= rack(0);
      type_cast_739_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_739_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp610x_xop_736,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_102_740,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_73_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_73_inst_req_0;
      type_cast_73_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_73_inst_req_1;
      type_cast_73_inst_ack_1<= rack(0);
      type_cast_73_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_73_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call13_67,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv18_74,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_762_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_762_inst_req_0;
      type_cast_762_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_762_inst_req_1;
      type_cast_762_inst_ack_1<= rack(0);
      type_cast_762_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_762_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext602_937,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_762_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_779_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_779_inst_req_0;
      type_cast_779_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_779_inst_req_1;
      type_cast_779_inst_ack_1<= rack(0);
      type_cast_779_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_779_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call313_773,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv316_780,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_795_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_795_inst_req_0;
      type_cast_795_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_795_inst_req_1;
      type_cast_795_inst_ack_1<= rack(0);
      type_cast_795_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_795_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call321_789,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv325_796,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_816_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_816_inst_req_0;
      type_cast_816_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_816_inst_req_1;
      type_cast_816_inst_ack_1<= rack(0);
      type_cast_816_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_816_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call331_810,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv335_817,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_837_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_837_inst_req_0;
      type_cast_837_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_837_inst_req_1;
      type_cast_837_inst_ack_1<= rack(0);
      type_cast_837_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_837_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call341_831,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv345_838,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_858_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_858_inst_req_0;
      type_cast_858_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_858_inst_req_1;
      type_cast_858_inst_ack_1<= rack(0);
      type_cast_858_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_858_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call351_852,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv355_859,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_879_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_879_inst_req_0;
      type_cast_879_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_879_inst_req_1;
      type_cast_879_inst_ack_1<= rack(0);
      type_cast_879_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_879_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call361_873,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv365_880,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_89_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_89_inst_req_0;
      type_cast_89_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_89_inst_req_1;
      type_cast_89_inst_ack_1<= rack(0);
      type_cast_89_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_89_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_83,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv25_90,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_900_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_900_inst_req_0;
      type_cast_900_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_900_inst_req_1;
      type_cast_900_inst_ack_1<= rack(0);
      type_cast_900_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_900_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call371_894,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv375_901,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_921_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_921_inst_req_0;
      type_cast_921_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_921_inst_req_1;
      type_cast_921_inst_ack_1<= rack(0);
      type_cast_921_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_921_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call381_915,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv385_922,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_954_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_954_inst_req_0;
      type_cast_954_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_954_inst_req_1;
      type_cast_954_inst_ack_1<= rack(0);
      type_cast_954_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_954_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add182_396,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv397_955,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_958_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_958_inst_req_0;
      type_cast_958_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_958_inst_req_1;
      type_cast_958_inst_ack_1<= rack(0);
      type_cast_958_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_958_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add199_427,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv399_959,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_962_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_962_inst_req_0;
      type_cast_962_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_962_inst_req_1;
      type_cast_962_inst_ack_1<= rack(0);
      type_cast_962_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_962_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add216_458,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv402_963,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1036_index_1_rename
    process(R_indvar587_1035_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar587_1035_resized;
      ov(13 downto 0) := iv;
      R_indvar587_1035_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1036_index_1_resize
    process(indvar587_1024) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar587_1024;
      ov := iv(13 downto 0);
      R_indvar587_1035_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1036_root_address_inst
    process(array_obj_ref_1036_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1036_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1036_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1302_index_1_rename
    process(R_indvar_1301_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1301_resized;
      ov(13 downto 0) := iv;
      R_indvar_1301_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1302_index_1_resize
    process(indvar_1290) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1290;
      ov := iv(13 downto 0);
      R_indvar_1301_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1302_root_address_inst
    process(array_obj_ref_1302_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1302_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1302_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_537_index_1_rename
    process(R_indvar617_536_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar617_536_resized;
      ov(13 downto 0) := iv;
      R_indvar617_536_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_537_index_1_resize
    process(indvar617_525) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar617_525;
      ov := iv(13 downto 0);
      R_indvar617_536_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_537_root_address_inst
    process(array_obj_ref_537_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_537_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_537_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_768_index_1_rename
    process(R_indvar601_767_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar601_767_resized;
      ov(10 downto 0) := iv;
      R_indvar601_767_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_768_index_1_resize
    process(indvar601_756) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar601_756;
      ov := iv(10 downto 0);
      R_indvar601_767_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_768_root_address_inst
    process(array_obj_ref_768_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_768_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_768_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1040_addr_0
    process(ptr_deref_1040_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1040_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1040_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1040_base_resize
    process(arrayidx413_1038) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx413_1038;
      ov := iv(13 downto 0);
      ptr_deref_1040_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1040_gather_scatter
    process(type_cast_1042_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1042_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1040_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1040_root_address_inst
    process(ptr_deref_1040_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1040_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1040_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1307_addr_0
    process(ptr_deref_1307_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1307_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1307_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1307_base_resize
    process(arrayidx495_1304) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx495_1304;
      ov := iv(13 downto 0);
      ptr_deref_1307_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1307_gather_scatter
    process(ptr_deref_1307_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1307_data_0;
      ov(63 downto 0) := iv;
      tmp496_1308 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1307_root_address_inst
    process(ptr_deref_1307_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1307_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1307_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_698_addr_0
    process(ptr_deref_698_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_698_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_698_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_698_base_resize
    process(arrayidx_539) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_539;
      ov := iv(13 downto 0);
      ptr_deref_698_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_698_gather_scatter
    process(add298_696) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add298_696;
      ov(63 downto 0) := iv;
      ptr_deref_698_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_698_root_address_inst
    process(ptr_deref_698_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_698_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_698_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_929_addr_0
    process(ptr_deref_929_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_929_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_929_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_929_base_resize
    process(arrayidx390_770) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx390_770;
      ov := iv(10 downto 0);
      ptr_deref_929_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_929_gather_scatter
    process(add386_927) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add386_927;
      ov(63 downto 0) := iv;
      ptr_deref_929_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_929_root_address_inst
    process(ptr_deref_929_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_929_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_929_root_address <= ov(10 downto 0);
      --
    end process;
    if_stmt_1055_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_1054;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1055_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1055_branch_req_0,
          ack0 => if_stmt_1055_branch_ack_0,
          ack1 => if_stmt_1055_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1246_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp408567_979;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1246_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1246_branch_req_0,
          ack0 => if_stmt_1246_branch_ack_0,
          ack1 => if_stmt_1246_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1418_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1417;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1418_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1418_branch_req_0,
          ack0 => if_stmt_1418_branch_ack_0,
          ack1 => if_stmt_1418_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_466_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp575_465;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_466_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_466_branch_req_0,
          ack0 => if_stmt_466_branch_ack_0,
          ack1 => if_stmt_466_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_481_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp306571_480;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_481_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_481_branch_req_0,
          ack0 => if_stmt_481_branch_ack_0,
          ack1 => if_stmt_481_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_712_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_711;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_712_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_712_branch_req_0,
          ack0 => if_stmt_712_branch_ack_0,
          ack1 => if_stmt_712_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_943_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_942;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_943_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_943_branch_req_0,
          ack0 => if_stmt_943_branch_ack_0,
          ack1 => if_stmt_943_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_980_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp408567_979;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_980_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_980_branch_req_0,
          ack0 => if_stmt_980_branch_ack_0,
          ack1 => if_stmt_980_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1003_inst
    process(tmp594_992) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp594_992, type_cast_1002_wire_constant, tmp_var);
      tmp594x_xop_1004 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1269_inst
    process(tmp582_1258) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp582_1258, type_cast_1268_wire_constant, tmp_var);
      tmp582x_xop_1270 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_504_inst
    process(tmp624_493) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp624_493, type_cast_503_wire_constant, tmp_var);
      tmp624x_xop_505 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_735_inst
    process(tmp610_724) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp610_724, type_cast_734_wire_constant, tmp_var);
      tmp610x_xop_736 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1013_inst
    process(iNsTr_132_1008) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_132_1008, type_cast_1012_wire_constant, tmp_var);
      xx_xop631_1014 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1048_inst
    process(indvar587_1024) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar587_1024, type_cast_1047_wire_constant, tmp_var);
      indvarx_xnext588_1049 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1279_inst
    process(iNsTr_243_1274) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_243_1274, type_cast_1278_wire_constant, tmp_var);
      xx_xop_1280 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1411_inst
    process(indvar_1290) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1290, type_cast_1410_wire_constant, tmp_var);
      indvarx_xnext_1412 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_514_inst
    process(iNsTr_73_509) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_73_509, type_cast_513_wire_constant, tmp_var);
      xx_xop633_515 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_705_inst
    process(indvar617_525) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar617_525, type_cast_704_wire_constant, tmp_var);
      indvarx_xnext618_706 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_745_inst
    process(iNsTr_102_740) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_102_740, type_cast_744_wire_constant, tmp_var);
      xx_xop632_746 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_936_inst
    process(indvar601_756) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar601_756, type_cast_935_wire_constant, tmp_var);
      indvarx_xnext602_937 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1053_inst
    process(indvarx_xnext588_1049, tmp599_1021) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext588_1049, tmp599_1021, tmp_var);
      exitcond_1054 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1416_inst
    process(indvarx_xnext_1412, tmp586_1287) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1412, tmp586_1287, tmp_var);
      exitcond1_1417 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_710_inst
    process(indvarx_xnext618_706, tmp629_522) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext618_706, tmp629_522, tmp_var);
      exitcond3_711 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_941_inst
    process(indvarx_xnext602_937, tmp615_753) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext602_937, tmp615_753, tmp_var);
      exitcond2_942 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1257_inst
    process(mul403_973) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul403_973, type_cast_1256_wire_constant, tmp_var);
      tmp582_1258 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_492_inst
    process(mul120_272) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul120_272, type_cast_491_wire_constant, tmp_var);
      tmp624_493 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_723_inst
    process(mul132_303) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul132_303, type_cast_722_wire_constant, tmp_var);
      tmp610_724 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_991_inst
    process(mul403_973) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul403_973, type_cast_990_wire_constant, tmp_var);
      tmp594_992 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1317_inst
    process(tmp496_1308) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp496_1308, type_cast_1316_wire_constant, tmp_var);
      shr502_1318 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1327_inst
    process(tmp496_1308) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp496_1308, type_cast_1326_wire_constant, tmp_var);
      shr508_1328 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1337_inst
    process(tmp496_1308) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp496_1308, type_cast_1336_wire_constant, tmp_var);
      shr514_1338 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1347_inst
    process(tmp496_1308) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp496_1308, type_cast_1346_wire_constant, tmp_var);
      shr520_1348 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1357_inst
    process(tmp496_1308) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp496_1308, type_cast_1356_wire_constant, tmp_var);
      shr526_1358 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1367_inst
    process(tmp496_1308) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp496_1308, type_cast_1366_wire_constant, tmp_var);
      shr532_1368 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1377_inst
    process(tmp496_1308) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp496_1308, type_cast_1376_wire_constant, tmp_var);
      shr538_1378 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_266_inst
    process(conv117_258, conv115_254) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv117_258, conv115_254, tmp_var);
      mul_267 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_271_inst
    process(mul_267, conv119_262) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_267, conv119_262, tmp_var);
      mul120_272 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_292_inst
    process(conv125_280, conv123_276) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv125_280, conv123_276, tmp_var);
      mul126_293 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_297_inst
    process(mul126_293, conv128_284) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul126_293, conv128_284, tmp_var);
      mul129_298 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_302_inst
    process(mul129_298, conv131_288) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul129_298, conv131_288, tmp_var);
      mul132_303 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_967_inst
    process(conv399_959, conv397_955) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv399_959, conv397_955, tmp_var);
      mul400_968 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_972_inst
    process(mul400_968, conv402_963) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul400_968, conv402_963, tmp_var);
      mul403_973 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_125_inst
    process(conv42_121, shl36_111) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv42_121, shl36_111, tmp_var);
      add43_126 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_156_inst
    process(conv59_152, shl53_142) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv59_152, shl53_142, tmp_var);
      add60_157 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_187_inst
    process(conv76_183, shl70_173) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv76_183, shl70_173, tmp_var);
      add77_188 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_218_inst
    process(conv93_214, shl87_204) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv93_214, shl87_204, tmp_var);
      add94_219 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_249_inst
    process(conv110_245, shl104_235) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv110_245, shl104_235, tmp_var);
      add111_250 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_333_inst
    process(conv147_329, shl141_319) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv147_329, shl141_319, tmp_var);
      add148_334 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_364_inst
    process(conv164_360, shl158_350) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv164_360, shl158_350, tmp_var);
      add165_365 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_395_inst
    process(conv181_391, shl175_381) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv181_391, shl175_381, tmp_var);
      add182_396 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_426_inst
    process(conv198_422, shl192_412) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv198_422, shl192_412, tmp_var);
      add199_427 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_457_inst
    process(conv215_453, shl209_443) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv215_453, shl209_443, tmp_var);
      add216_458 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_63_inst
    process(conv9_59, shl_49) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv9_59, shl_49, tmp_var);
      add_64 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_94_inst
    process(conv25_90, shl19_80) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv25_90, shl19_80, tmp_var);
      add26_95 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_569_inst
    process(conv237_565, shl230_555) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv237_565, shl230_555, tmp_var);
      add238_570 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_590_inst
    process(shl240_576, conv247_586) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl240_576, conv247_586, tmp_var);
      add248_591 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_611_inst
    process(shl250_597, conv257_607) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl250_597, conv257_607, tmp_var);
      add258_612 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_632_inst
    process(shl260_618, conv267_628) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl260_618, conv267_628, tmp_var);
      add268_633 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_653_inst
    process(shl270_639, conv277_649) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl270_639, conv277_649, tmp_var);
      add278_654 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_674_inst
    process(shl280_660, conv287_670) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl280_660, conv287_670, tmp_var);
      add288_675 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_695_inst
    process(shl290_681, conv297_691) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl290_681, conv297_691, tmp_var);
      add298_696 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_800_inst
    process(conv325_796, shl318_786) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv325_796, shl318_786, tmp_var);
      add326_801 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_821_inst
    process(shl328_807, conv335_817) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl328_807, conv335_817, tmp_var);
      add336_822 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_842_inst
    process(shl338_828, conv345_838) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl338_828, conv345_838, tmp_var);
      add346_843 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_863_inst
    process(shl348_849, conv355_859) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl348_849, conv355_859, tmp_var);
      add356_864 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_884_inst
    process(shl358_870, conv365_880) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl358_870, conv365_880, tmp_var);
      add366_885 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_905_inst
    process(shl368_891, conv375_901) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl368_891, conv375_901, tmp_var);
      add376_906 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_926_inst
    process(shl378_912, conv385_922) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl378_912, conv385_922, tmp_var);
      add386_927 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_110_inst
    process(conv35_105) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_105, type_cast_109_wire_constant, tmp_var);
      shl36_111 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_141_inst
    process(conv52_136) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv52_136, type_cast_140_wire_constant, tmp_var);
      shl53_142 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_172_inst
    process(conv69_167) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv69_167, type_cast_171_wire_constant, tmp_var);
      shl70_173 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_203_inst
    process(conv86_198) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv86_198, type_cast_202_wire_constant, tmp_var);
      shl87_204 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_234_inst
    process(conv103_229) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv103_229, type_cast_233_wire_constant, tmp_var);
      shl104_235 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_318_inst
    process(conv140_313) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv140_313, type_cast_317_wire_constant, tmp_var);
      shl141_319 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_349_inst
    process(conv157_344) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv157_344, type_cast_348_wire_constant, tmp_var);
      shl158_350 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_380_inst
    process(conv174_375) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv174_375, type_cast_379_wire_constant, tmp_var);
      shl175_381 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_411_inst
    process(conv191_406) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv191_406, type_cast_410_wire_constant, tmp_var);
      shl192_412 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_442_inst
    process(conv208_437) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv208_437, type_cast_441_wire_constant, tmp_var);
      shl209_443 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_48_inst
    process(conv3_43) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv3_43, type_cast_47_wire_constant, tmp_var);
      shl_49 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_79_inst
    process(conv18_74) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv18_74, type_cast_78_wire_constant, tmp_var);
      shl19_80 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_554_inst
    process(conv228_549) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv228_549, type_cast_553_wire_constant, tmp_var);
      shl230_555 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_575_inst
    process(add238_570) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add238_570, type_cast_574_wire_constant, tmp_var);
      shl240_576 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_596_inst
    process(add248_591) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add248_591, type_cast_595_wire_constant, tmp_var);
      shl250_597 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_617_inst
    process(add258_612) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add258_612, type_cast_616_wire_constant, tmp_var);
      shl260_618 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_638_inst
    process(add268_633) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add268_633, type_cast_637_wire_constant, tmp_var);
      shl270_639 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_659_inst
    process(add278_654) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add278_654, type_cast_658_wire_constant, tmp_var);
      shl280_660 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_680_inst
    process(add288_675) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add288_675, type_cast_679_wire_constant, tmp_var);
      shl290_681 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_785_inst
    process(conv316_780) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv316_780, type_cast_784_wire_constant, tmp_var);
      shl318_786 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_806_inst
    process(add326_801) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add326_801, type_cast_805_wire_constant, tmp_var);
      shl328_807 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_827_inst
    process(add336_822) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add336_822, type_cast_826_wire_constant, tmp_var);
      shl338_828 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_848_inst
    process(add346_843) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add346_843, type_cast_847_wire_constant, tmp_var);
      shl348_849 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_869_inst
    process(add356_864) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add356_864, type_cast_868_wire_constant, tmp_var);
      shl358_870 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_890_inst
    process(add366_885) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add366_885, type_cast_889_wire_constant, tmp_var);
      shl368_891 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_911_inst
    process(add376_906) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add376_906, type_cast_910_wire_constant, tmp_var);
      shl378_912 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1240_inst
    process(conv479_1236, conv420_1072) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv479_1236, conv420_1072, tmp_var);
      sub_1241 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1263_inst
    process(tmp582_1258) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp582_1258, type_cast_1262_wire_constant, tmp_var);
      tmp583_1264 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_463_inst
    process(mul120_272) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul120_272, type_cast_462_wire_constant, tmp_var);
      cmp575_465 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_479_inst
    process(mul132_303) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul132_303, type_cast_478_wire_constant, tmp_var);
      cmp306571_480 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_498_inst
    process(tmp624_493) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp624_493, type_cast_497_wire_constant, tmp_var);
      tmp625_499 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_729_inst
    process(tmp610_724) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp610_724, type_cast_728_wire_constant, tmp_var);
      tmp611_730 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_978_inst
    process(mul403_973) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul403_973, type_cast_977_wire_constant, tmp_var);
      cmp408567_979 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_997_inst
    process(tmp594_992) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp594_992, type_cast_996_wire_constant, tmp_var);
      tmp595_998 <= tmp_var; --
    end process;
    -- shared split operator group (94) : array_obj_ref_1036_index_offset 
    ApIntAdd_group_94: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar587_1035_scaled;
      array_obj_ref_1036_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1036_index_offset_req_0;
      array_obj_ref_1036_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1036_index_offset_req_1;
      array_obj_ref_1036_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_94_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_94_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_94",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 94
    -- shared split operator group (95) : array_obj_ref_1302_index_offset 
    ApIntAdd_group_95: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1301_scaled;
      array_obj_ref_1302_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1302_index_offset_req_0;
      array_obj_ref_1302_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1302_index_offset_req_1;
      array_obj_ref_1302_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_95_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_95_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_95",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 95
    -- shared split operator group (96) : array_obj_ref_537_index_offset 
    ApIntAdd_group_96: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar617_536_scaled;
      array_obj_ref_537_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_537_index_offset_req_0;
      array_obj_ref_537_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_537_index_offset_req_1;
      array_obj_ref_537_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_96_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_96_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_96",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 96
    -- shared split operator group (97) : array_obj_ref_768_index_offset 
    ApIntAdd_group_97: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar601_767_scaled;
      array_obj_ref_768_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_768_index_offset_req_0;
      array_obj_ref_768_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_768_index_offset_req_1;
      array_obj_ref_768_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_97_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_97_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_97",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100010",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 97
    -- unary operator type_cast_1070_inst
    process(call419_1066) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call419_1066, tmp_var);
      type_cast_1070_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1234_inst
    process(call478_1231) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call478_1231, tmp_var);
      type_cast_1234_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1307_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1307_load_0_req_0;
      ptr_deref_1307_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1307_load_0_req_1;
      ptr_deref_1307_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1307_word_address_0;
      ptr_deref_1307_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1040_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1040_store_0_req_0;
      ptr_deref_1040_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1040_store_0_req_1;
      ptr_deref_1040_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1040_word_address_0;
      data_in <= ptr_deref_1040_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_698_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_698_store_0_req_0;
      ptr_deref_698_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_698_store_0_req_1;
      ptr_deref_698_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_698_word_address_0;
      data_in <= ptr_deref_698_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_929_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_929_store_0_req_0;
      ptr_deref_929_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_929_store_0_req_1;
      ptr_deref_929_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_929_word_address_0;
      data_in <= ptr_deref_929_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(10 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_Block0_done_1218_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1218_inst_req_0;
      RPIPE_Block0_done_1218_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1218_inst_req_1;
      RPIPE_Block0_done_1218_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call470_1219 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1221_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1221_inst_req_0;
      RPIPE_Block1_done_1221_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1221_inst_req_1;
      RPIPE_Block1_done_1221_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call472_1222 <= data_out(15 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1224_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1224_inst_req_0;
      RPIPE_Block2_done_1224_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1224_inst_req_1;
      RPIPE_Block2_done_1224_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call474_1225 <= data_out(15 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1227_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1227_inst_req_0;
      RPIPE_Block3_done_1227_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1227_inst_req_1;
      RPIPE_Block3_done_1227_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call476_1228 <= data_out(15 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_ConvTranspose_input_pipe_599_inst RPIPE_ConvTranspose_input_pipe_683_inst RPIPE_ConvTranspose_input_pipe_788_inst RPIPE_ConvTranspose_input_pipe_541_inst RPIPE_ConvTranspose_input_pipe_578_inst RPIPE_ConvTranspose_input_pipe_772_inst RPIPE_ConvTranspose_input_pipe_620_inst RPIPE_ConvTranspose_input_pipe_35_inst RPIPE_ConvTranspose_input_pipe_641_inst RPIPE_ConvTranspose_input_pipe_557_inst RPIPE_ConvTranspose_input_pipe_662_inst RPIPE_ConvTranspose_input_pipe_809_inst RPIPE_ConvTranspose_input_pipe_872_inst RPIPE_ConvTranspose_input_pipe_830_inst RPIPE_ConvTranspose_input_pipe_851_inst RPIPE_ConvTranspose_input_pipe_893_inst RPIPE_ConvTranspose_input_pipe_914_inst RPIPE_ConvTranspose_input_pipe_51_inst RPIPE_ConvTranspose_input_pipe_66_inst RPIPE_ConvTranspose_input_pipe_82_inst RPIPE_ConvTranspose_input_pipe_97_inst RPIPE_ConvTranspose_input_pipe_113_inst RPIPE_ConvTranspose_input_pipe_128_inst RPIPE_ConvTranspose_input_pipe_144_inst RPIPE_ConvTranspose_input_pipe_159_inst RPIPE_ConvTranspose_input_pipe_175_inst RPIPE_ConvTranspose_input_pipe_190_inst RPIPE_ConvTranspose_input_pipe_206_inst RPIPE_ConvTranspose_input_pipe_221_inst RPIPE_ConvTranspose_input_pipe_237_inst RPIPE_ConvTranspose_input_pipe_305_inst RPIPE_ConvTranspose_input_pipe_321_inst RPIPE_ConvTranspose_input_pipe_336_inst RPIPE_ConvTranspose_input_pipe_352_inst RPIPE_ConvTranspose_input_pipe_367_inst RPIPE_ConvTranspose_input_pipe_383_inst RPIPE_ConvTranspose_input_pipe_398_inst RPIPE_ConvTranspose_input_pipe_414_inst RPIPE_ConvTranspose_input_pipe_429_inst RPIPE_ConvTranspose_input_pipe_445_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(319 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 39 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 39 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 39 downto 0);
      signal guard_vector : std_logic_vector( 39 downto 0);
      constant outBUFs : IntegerArray(39 downto 0) := (39 => 1, 38 => 1, 37 => 1, 36 => 1, 35 => 1, 34 => 1, 33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(39 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false, 35 => false, 36 => false, 37 => false, 38 => false, 39 => false);
      constant guardBuffering: IntegerArray(39 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2, 35 => 2, 36 => 2, 37 => 2, 38 => 2, 39 => 2);
      -- 
    begin -- 
      reqL_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_599_inst_req_0;
      reqL_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_683_inst_req_0;
      reqL_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_788_inst_req_0;
      reqL_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_541_inst_req_0;
      reqL_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_578_inst_req_0;
      reqL_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_772_inst_req_0;
      reqL_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_620_inst_req_0;
      reqL_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_35_inst_req_0;
      reqL_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_641_inst_req_0;
      reqL_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_557_inst_req_0;
      reqL_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_662_inst_req_0;
      reqL_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_809_inst_req_0;
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_872_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_830_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_851_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_893_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_914_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_51_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_66_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_82_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_97_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_113_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_128_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_144_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_159_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_175_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_190_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_206_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_221_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_237_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_305_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_321_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_336_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_352_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_367_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_383_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_398_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_414_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_429_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_445_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_599_inst_ack_0 <= ackL_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_683_inst_ack_0 <= ackL_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_788_inst_ack_0 <= ackL_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_541_inst_ack_0 <= ackL_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_578_inst_ack_0 <= ackL_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_772_inst_ack_0 <= ackL_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_620_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_35_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_641_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_557_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_662_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_809_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_872_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_830_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_851_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_893_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_914_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_51_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_66_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_82_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_97_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_113_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_128_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_144_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_159_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_175_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_190_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_206_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_221_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_237_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_305_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_321_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_336_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_352_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_367_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_383_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_398_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_414_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_429_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_445_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_599_inst_req_1;
      reqR_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_683_inst_req_1;
      reqR_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_788_inst_req_1;
      reqR_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_541_inst_req_1;
      reqR_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_578_inst_req_1;
      reqR_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_772_inst_req_1;
      reqR_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_620_inst_req_1;
      reqR_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_35_inst_req_1;
      reqR_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_641_inst_req_1;
      reqR_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_557_inst_req_1;
      reqR_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_662_inst_req_1;
      reqR_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_809_inst_req_1;
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_872_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_830_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_851_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_893_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_914_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_51_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_66_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_82_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_97_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_113_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_128_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_144_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_159_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_175_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_190_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_206_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_221_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_237_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_305_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_321_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_336_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_352_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_367_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_383_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_398_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_414_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_429_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_445_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_599_inst_ack_1 <= ackR_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_683_inst_ack_1 <= ackR_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_788_inst_ack_1 <= ackR_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_541_inst_ack_1 <= ackR_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_578_inst_ack_1 <= ackR_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_772_inst_ack_1 <= ackR_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_620_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_35_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_641_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_557_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_662_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_809_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_872_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_830_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_851_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_893_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_914_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_51_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_66_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_82_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_97_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_113_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_128_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_144_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_159_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_175_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_190_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_206_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_221_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_237_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_305_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_321_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_336_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_352_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_367_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_383_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_398_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_414_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_429_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_445_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      call253_600 <= data_out(319 downto 312);
      call293_684 <= data_out(311 downto 304);
      call321_789 <= data_out(303 downto 296);
      call225_542 <= data_out(295 downto 288);
      call243_579 <= data_out(287 downto 280);
      call313_773 <= data_out(279 downto 272);
      call263_621 <= data_out(271 downto 264);
      call_36 <= data_out(263 downto 256);
      call273_642 <= data_out(255 downto 248);
      call233_558 <= data_out(247 downto 240);
      call283_663 <= data_out(239 downto 232);
      call331_810 <= data_out(231 downto 224);
      call361_873 <= data_out(223 downto 216);
      call341_831 <= data_out(215 downto 208);
      call351_852 <= data_out(207 downto 200);
      call371_894 <= data_out(199 downto 192);
      call381_915 <= data_out(191 downto 184);
      call6_52 <= data_out(183 downto 176);
      call13_67 <= data_out(175 downto 168);
      call22_83 <= data_out(167 downto 160);
      call30_98 <= data_out(159 downto 152);
      call39_114 <= data_out(151 downto 144);
      call47_129 <= data_out(143 downto 136);
      call56_145 <= data_out(135 downto 128);
      call64_160 <= data_out(127 downto 120);
      call73_176 <= data_out(119 downto 112);
      call81_191 <= data_out(111 downto 104);
      call90_207 <= data_out(103 downto 96);
      call98_222 <= data_out(95 downto 88);
      call107_238 <= data_out(87 downto 80);
      call135_306 <= data_out(79 downto 72);
      call144_322 <= data_out(71 downto 64);
      call152_337 <= data_out(63 downto 56);
      call161_353 <= data_out(55 downto 48);
      call169_368 <= data_out(47 downto 40);
      call178_384 <= data_out(39 downto 32);
      call186_399 <= data_out(31 downto 24);
      call195_415 <= data_out(23 downto 16);
      call203_430 <= data_out(15 downto 8);
      call212_446 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_4_gI", nreqs => 40, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_4: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_4", data_width => 8,  num_reqs => 40,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared outport operator group (0) : WPIPE_Block0_start_1073_inst WPIPE_Block0_start_1076_inst WPIPE_Block0_start_1079_inst WPIPE_Block0_start_1082_inst WPIPE_Block0_start_1085_inst WPIPE_Block0_start_1088_inst WPIPE_Block0_start_1091_inst WPIPE_Block0_start_1094_inst WPIPE_Block0_start_1097_inst WPIPE_Block0_start_1100_inst WPIPE_Block0_start_1103_inst WPIPE_Block0_start_1106_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal sample_req, sample_ack : BooleanArray( 11 downto 0);
      signal update_req, update_ack : BooleanArray( 11 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 11 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant inBUFs : IntegerArray(11 downto 0) := (11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      sample_req_unguarded(11) <= WPIPE_Block0_start_1073_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block0_start_1076_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block0_start_1079_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block0_start_1082_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block0_start_1085_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block0_start_1088_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block0_start_1091_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block0_start_1094_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block0_start_1097_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block0_start_1100_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block0_start_1103_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block0_start_1106_inst_req_0;
      WPIPE_Block0_start_1073_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block0_start_1076_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block0_start_1079_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block0_start_1082_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block0_start_1085_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block0_start_1088_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block0_start_1091_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block0_start_1094_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block0_start_1097_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block0_start_1100_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block0_start_1103_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block0_start_1106_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(11) <= WPIPE_Block0_start_1073_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block0_start_1076_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block0_start_1079_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block0_start_1082_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block0_start_1085_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block0_start_1088_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block0_start_1091_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block0_start_1094_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block0_start_1097_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block0_start_1100_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block0_start_1103_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block0_start_1106_inst_req_1;
      WPIPE_Block0_start_1073_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block0_start_1076_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block0_start_1079_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block0_start_1082_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block0_start_1085_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block0_start_1088_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block0_start_1091_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block0_start_1094_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block0_start_1097_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block0_start_1100_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block0_start_1103_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block0_start_1106_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      data_in <= add_64 & add26_95 & add43_126 & add60_157 & add77_188 & add94_219 & add111_250 & add148_334 & add165_365 & add182_396 & add199_427 & add216_458;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 12, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_1112_inst WPIPE_Block1_start_1142_inst WPIPE_Block1_start_1130_inst WPIPE_Block1_start_1121_inst WPIPE_Block1_start_1139_inst WPIPE_Block1_start_1109_inst WPIPE_Block1_start_1133_inst WPIPE_Block1_start_1127_inst WPIPE_Block1_start_1115_inst WPIPE_Block1_start_1124_inst WPIPE_Block1_start_1136_inst WPIPE_Block1_start_1118_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal sample_req, sample_ack : BooleanArray( 11 downto 0);
      signal update_req, update_ack : BooleanArray( 11 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 11 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant inBUFs : IntegerArray(11 downto 0) := (11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      sample_req_unguarded(11) <= WPIPE_Block1_start_1112_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block1_start_1142_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block1_start_1130_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block1_start_1121_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block1_start_1139_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block1_start_1109_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block1_start_1133_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block1_start_1127_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block1_start_1115_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block1_start_1124_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block1_start_1136_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block1_start_1118_inst_req_0;
      WPIPE_Block1_start_1112_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block1_start_1142_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block1_start_1130_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block1_start_1121_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block1_start_1139_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block1_start_1109_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block1_start_1133_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block1_start_1127_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block1_start_1115_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block1_start_1124_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block1_start_1136_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block1_start_1118_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(11) <= WPIPE_Block1_start_1112_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block1_start_1142_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block1_start_1130_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block1_start_1121_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block1_start_1139_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block1_start_1109_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block1_start_1133_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block1_start_1127_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block1_start_1115_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block1_start_1124_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block1_start_1136_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block1_start_1118_inst_req_1;
      WPIPE_Block1_start_1112_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block1_start_1142_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block1_start_1130_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block1_start_1121_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block1_start_1139_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block1_start_1109_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block1_start_1133_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block1_start_1127_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block1_start_1115_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block1_start_1124_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block1_start_1136_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block1_start_1118_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      data_in <= add26_95 & add216_458 & add148_334 & add77_188 & add199_427 & add_64 & add165_365 & add111_250 & add43_126 & add94_219 & add182_396 & add60_157;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 16, num_reqs => 12, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1145_inst WPIPE_Block2_start_1157_inst WPIPE_Block2_start_1151_inst WPIPE_Block2_start_1160_inst WPIPE_Block2_start_1172_inst WPIPE_Block2_start_1148_inst WPIPE_Block2_start_1175_inst WPIPE_Block2_start_1154_inst WPIPE_Block2_start_1166_inst WPIPE_Block2_start_1178_inst WPIPE_Block2_start_1163_inst WPIPE_Block2_start_1169_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal sample_req, sample_ack : BooleanArray( 11 downto 0);
      signal update_req, update_ack : BooleanArray( 11 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 11 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant inBUFs : IntegerArray(11 downto 0) := (11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      sample_req_unguarded(11) <= WPIPE_Block2_start_1145_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block2_start_1157_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block2_start_1151_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block2_start_1160_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block2_start_1172_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block2_start_1148_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block2_start_1175_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block2_start_1154_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block2_start_1166_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block2_start_1178_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block2_start_1163_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block2_start_1169_inst_req_0;
      WPIPE_Block2_start_1145_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block2_start_1157_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block2_start_1151_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block2_start_1160_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block2_start_1172_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block2_start_1148_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block2_start_1175_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block2_start_1154_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block2_start_1166_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block2_start_1178_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block2_start_1163_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block2_start_1169_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(11) <= WPIPE_Block2_start_1145_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block2_start_1157_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block2_start_1151_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block2_start_1160_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block2_start_1172_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block2_start_1148_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block2_start_1175_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block2_start_1154_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block2_start_1166_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block2_start_1178_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block2_start_1163_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block2_start_1169_inst_req_1;
      WPIPE_Block2_start_1145_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block2_start_1157_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block2_start_1151_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block2_start_1160_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block2_start_1172_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block2_start_1148_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block2_start_1175_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block2_start_1154_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block2_start_1166_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block2_start_1178_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block2_start_1163_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block2_start_1169_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      data_in <= add_64 & add77_188 & add43_126 & add94_219 & add182_396 & add26_95 & add199_427 & add60_157 & add148_334 & add216_458 & add111_250 & add165_365;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 16, num_reqs => 12, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1181_inst WPIPE_Block3_start_1184_inst WPIPE_Block3_start_1187_inst WPIPE_Block3_start_1190_inst WPIPE_Block3_start_1196_inst WPIPE_Block3_start_1193_inst WPIPE_Block3_start_1211_inst WPIPE_Block3_start_1205_inst WPIPE_Block3_start_1199_inst WPIPE_Block3_start_1214_inst WPIPE_Block3_start_1208_inst WPIPE_Block3_start_1202_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal sample_req, sample_ack : BooleanArray( 11 downto 0);
      signal update_req, update_ack : BooleanArray( 11 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 11 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant inBUFs : IntegerArray(11 downto 0) := (11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      sample_req_unguarded(11) <= WPIPE_Block3_start_1181_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block3_start_1184_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block3_start_1187_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block3_start_1190_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block3_start_1196_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block3_start_1193_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block3_start_1211_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block3_start_1205_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block3_start_1199_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block3_start_1214_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block3_start_1208_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block3_start_1202_inst_req_0;
      WPIPE_Block3_start_1181_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block3_start_1184_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block3_start_1187_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block3_start_1190_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block3_start_1196_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block3_start_1193_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block3_start_1211_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block3_start_1205_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block3_start_1199_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block3_start_1214_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block3_start_1208_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block3_start_1202_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(11) <= WPIPE_Block3_start_1181_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block3_start_1184_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block3_start_1187_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block3_start_1190_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block3_start_1196_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block3_start_1193_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block3_start_1211_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block3_start_1205_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block3_start_1199_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block3_start_1214_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block3_start_1208_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block3_start_1202_inst_req_1;
      WPIPE_Block3_start_1181_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block3_start_1184_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block3_start_1187_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block3_start_1190_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block3_start_1196_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block3_start_1193_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block3_start_1211_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block3_start_1205_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block3_start_1199_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block3_start_1214_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block3_start_1208_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block3_start_1202_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      data_in <= add_64 & add26_95 & add43_126 & add60_157 & add94_219 & add77_188 & add199_427 & add165_365 & add111_250 & add216_458 & add182_396 & add148_334;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 16, num_reqs => 12, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_ConvTranspose_output_pipe_790_inst WPIPE_ConvTranspose_output_pipe_580_inst WPIPE_ConvTranspose_output_pipe_774_inst WPIPE_ConvTranspose_output_pipe_543_inst WPIPE_ConvTranspose_output_pipe_601_inst WPIPE_ConvTranspose_output_pipe_685_inst WPIPE_ConvTranspose_output_pipe_622_inst WPIPE_ConvTranspose_output_pipe_37_inst WPIPE_ConvTranspose_output_pipe_643_inst WPIPE_ConvTranspose_output_pipe_664_inst WPIPE_ConvTranspose_output_pipe_874_inst WPIPE_ConvTranspose_output_pipe_811_inst WPIPE_ConvTranspose_output_pipe_559_inst WPIPE_ConvTranspose_output_pipe_832_inst WPIPE_ConvTranspose_output_pipe_853_inst WPIPE_ConvTranspose_output_pipe_895_inst WPIPE_ConvTranspose_output_pipe_916_inst WPIPE_ConvTranspose_output_pipe_53_inst WPIPE_ConvTranspose_output_pipe_68_inst WPIPE_ConvTranspose_output_pipe_84_inst WPIPE_ConvTranspose_output_pipe_99_inst WPIPE_ConvTranspose_output_pipe_115_inst WPIPE_ConvTranspose_output_pipe_130_inst WPIPE_ConvTranspose_output_pipe_146_inst WPIPE_ConvTranspose_output_pipe_161_inst WPIPE_ConvTranspose_output_pipe_177_inst WPIPE_ConvTranspose_output_pipe_192_inst WPIPE_ConvTranspose_output_pipe_208_inst WPIPE_ConvTranspose_output_pipe_223_inst WPIPE_ConvTranspose_output_pipe_239_inst WPIPE_ConvTranspose_output_pipe_307_inst WPIPE_ConvTranspose_output_pipe_323_inst WPIPE_ConvTranspose_output_pipe_338_inst WPIPE_ConvTranspose_output_pipe_354_inst WPIPE_ConvTranspose_output_pipe_369_inst WPIPE_ConvTranspose_output_pipe_385_inst WPIPE_ConvTranspose_output_pipe_400_inst WPIPE_ConvTranspose_output_pipe_416_inst WPIPE_ConvTranspose_output_pipe_431_inst WPIPE_ConvTranspose_output_pipe_447_inst WPIPE_ConvTranspose_output_pipe_1383_inst WPIPE_ConvTranspose_output_pipe_1386_inst WPIPE_ConvTranspose_output_pipe_1389_inst WPIPE_ConvTranspose_output_pipe_1392_inst WPIPE_ConvTranspose_output_pipe_1395_inst WPIPE_ConvTranspose_output_pipe_1398_inst WPIPE_ConvTranspose_output_pipe_1401_inst WPIPE_ConvTranspose_output_pipe_1404_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(383 downto 0);
      signal sample_req, sample_ack : BooleanArray( 47 downto 0);
      signal update_req, update_ack : BooleanArray( 47 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 47 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 47 downto 0);
      signal guard_vector : std_logic_vector( 47 downto 0);
      constant inBUFs : IntegerArray(47 downto 0) := (47 => 0, 46 => 0, 45 => 0, 44 => 0, 43 => 0, 42 => 0, 41 => 0, 40 => 0, 39 => 0, 38 => 0, 37 => 0, 36 => 0, 35 => 0, 34 => 0, 33 => 0, 32 => 0, 31 => 0, 30 => 0, 29 => 0, 28 => 0, 27 => 0, 26 => 0, 25 => 0, 24 => 0, 23 => 0, 22 => 0, 21 => 0, 20 => 0, 19 => 0, 18 => 0, 17 => 0, 16 => 0, 15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(47 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false, 35 => false, 36 => false, 37 => false, 38 => false, 39 => false, 40 => false, 41 => false, 42 => false, 43 => false, 44 => false, 45 => false, 46 => false, 47 => false);
      constant guardBuffering: IntegerArray(47 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2, 35 => 2, 36 => 2, 37 => 2, 38 => 2, 39 => 2, 40 => 2, 41 => 2, 42 => 2, 43 => 2, 44 => 2, 45 => 2, 46 => 2, 47 => 2);
      -- 
    begin -- 
      sample_req_unguarded(47) <= WPIPE_ConvTranspose_output_pipe_790_inst_req_0;
      sample_req_unguarded(46) <= WPIPE_ConvTranspose_output_pipe_580_inst_req_0;
      sample_req_unguarded(45) <= WPIPE_ConvTranspose_output_pipe_774_inst_req_0;
      sample_req_unguarded(44) <= WPIPE_ConvTranspose_output_pipe_543_inst_req_0;
      sample_req_unguarded(43) <= WPIPE_ConvTranspose_output_pipe_601_inst_req_0;
      sample_req_unguarded(42) <= WPIPE_ConvTranspose_output_pipe_685_inst_req_0;
      sample_req_unguarded(41) <= WPIPE_ConvTranspose_output_pipe_622_inst_req_0;
      sample_req_unguarded(40) <= WPIPE_ConvTranspose_output_pipe_37_inst_req_0;
      sample_req_unguarded(39) <= WPIPE_ConvTranspose_output_pipe_643_inst_req_0;
      sample_req_unguarded(38) <= WPIPE_ConvTranspose_output_pipe_664_inst_req_0;
      sample_req_unguarded(37) <= WPIPE_ConvTranspose_output_pipe_874_inst_req_0;
      sample_req_unguarded(36) <= WPIPE_ConvTranspose_output_pipe_811_inst_req_0;
      sample_req_unguarded(35) <= WPIPE_ConvTranspose_output_pipe_559_inst_req_0;
      sample_req_unguarded(34) <= WPIPE_ConvTranspose_output_pipe_832_inst_req_0;
      sample_req_unguarded(33) <= WPIPE_ConvTranspose_output_pipe_853_inst_req_0;
      sample_req_unguarded(32) <= WPIPE_ConvTranspose_output_pipe_895_inst_req_0;
      sample_req_unguarded(31) <= WPIPE_ConvTranspose_output_pipe_916_inst_req_0;
      sample_req_unguarded(30) <= WPIPE_ConvTranspose_output_pipe_53_inst_req_0;
      sample_req_unguarded(29) <= WPIPE_ConvTranspose_output_pipe_68_inst_req_0;
      sample_req_unguarded(28) <= WPIPE_ConvTranspose_output_pipe_84_inst_req_0;
      sample_req_unguarded(27) <= WPIPE_ConvTranspose_output_pipe_99_inst_req_0;
      sample_req_unguarded(26) <= WPIPE_ConvTranspose_output_pipe_115_inst_req_0;
      sample_req_unguarded(25) <= WPIPE_ConvTranspose_output_pipe_130_inst_req_0;
      sample_req_unguarded(24) <= WPIPE_ConvTranspose_output_pipe_146_inst_req_0;
      sample_req_unguarded(23) <= WPIPE_ConvTranspose_output_pipe_161_inst_req_0;
      sample_req_unguarded(22) <= WPIPE_ConvTranspose_output_pipe_177_inst_req_0;
      sample_req_unguarded(21) <= WPIPE_ConvTranspose_output_pipe_192_inst_req_0;
      sample_req_unguarded(20) <= WPIPE_ConvTranspose_output_pipe_208_inst_req_0;
      sample_req_unguarded(19) <= WPIPE_ConvTranspose_output_pipe_223_inst_req_0;
      sample_req_unguarded(18) <= WPIPE_ConvTranspose_output_pipe_239_inst_req_0;
      sample_req_unguarded(17) <= WPIPE_ConvTranspose_output_pipe_307_inst_req_0;
      sample_req_unguarded(16) <= WPIPE_ConvTranspose_output_pipe_323_inst_req_0;
      sample_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_338_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_354_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_369_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_385_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_400_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_416_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_431_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_447_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1383_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1386_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1389_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1392_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1395_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1398_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1401_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1404_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_790_inst_ack_0 <= sample_ack_unguarded(47);
      WPIPE_ConvTranspose_output_pipe_580_inst_ack_0 <= sample_ack_unguarded(46);
      WPIPE_ConvTranspose_output_pipe_774_inst_ack_0 <= sample_ack_unguarded(45);
      WPIPE_ConvTranspose_output_pipe_543_inst_ack_0 <= sample_ack_unguarded(44);
      WPIPE_ConvTranspose_output_pipe_601_inst_ack_0 <= sample_ack_unguarded(43);
      WPIPE_ConvTranspose_output_pipe_685_inst_ack_0 <= sample_ack_unguarded(42);
      WPIPE_ConvTranspose_output_pipe_622_inst_ack_0 <= sample_ack_unguarded(41);
      WPIPE_ConvTranspose_output_pipe_37_inst_ack_0 <= sample_ack_unguarded(40);
      WPIPE_ConvTranspose_output_pipe_643_inst_ack_0 <= sample_ack_unguarded(39);
      WPIPE_ConvTranspose_output_pipe_664_inst_ack_0 <= sample_ack_unguarded(38);
      WPIPE_ConvTranspose_output_pipe_874_inst_ack_0 <= sample_ack_unguarded(37);
      WPIPE_ConvTranspose_output_pipe_811_inst_ack_0 <= sample_ack_unguarded(36);
      WPIPE_ConvTranspose_output_pipe_559_inst_ack_0 <= sample_ack_unguarded(35);
      WPIPE_ConvTranspose_output_pipe_832_inst_ack_0 <= sample_ack_unguarded(34);
      WPIPE_ConvTranspose_output_pipe_853_inst_ack_0 <= sample_ack_unguarded(33);
      WPIPE_ConvTranspose_output_pipe_895_inst_ack_0 <= sample_ack_unguarded(32);
      WPIPE_ConvTranspose_output_pipe_916_inst_ack_0 <= sample_ack_unguarded(31);
      WPIPE_ConvTranspose_output_pipe_53_inst_ack_0 <= sample_ack_unguarded(30);
      WPIPE_ConvTranspose_output_pipe_68_inst_ack_0 <= sample_ack_unguarded(29);
      WPIPE_ConvTranspose_output_pipe_84_inst_ack_0 <= sample_ack_unguarded(28);
      WPIPE_ConvTranspose_output_pipe_99_inst_ack_0 <= sample_ack_unguarded(27);
      WPIPE_ConvTranspose_output_pipe_115_inst_ack_0 <= sample_ack_unguarded(26);
      WPIPE_ConvTranspose_output_pipe_130_inst_ack_0 <= sample_ack_unguarded(25);
      WPIPE_ConvTranspose_output_pipe_146_inst_ack_0 <= sample_ack_unguarded(24);
      WPIPE_ConvTranspose_output_pipe_161_inst_ack_0 <= sample_ack_unguarded(23);
      WPIPE_ConvTranspose_output_pipe_177_inst_ack_0 <= sample_ack_unguarded(22);
      WPIPE_ConvTranspose_output_pipe_192_inst_ack_0 <= sample_ack_unguarded(21);
      WPIPE_ConvTranspose_output_pipe_208_inst_ack_0 <= sample_ack_unguarded(20);
      WPIPE_ConvTranspose_output_pipe_223_inst_ack_0 <= sample_ack_unguarded(19);
      WPIPE_ConvTranspose_output_pipe_239_inst_ack_0 <= sample_ack_unguarded(18);
      WPIPE_ConvTranspose_output_pipe_307_inst_ack_0 <= sample_ack_unguarded(17);
      WPIPE_ConvTranspose_output_pipe_323_inst_ack_0 <= sample_ack_unguarded(16);
      WPIPE_ConvTranspose_output_pipe_338_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_354_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_369_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_385_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_400_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_416_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_431_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_447_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1383_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1386_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1389_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1392_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1395_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1398_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1401_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1404_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(47) <= WPIPE_ConvTranspose_output_pipe_790_inst_req_1;
      update_req_unguarded(46) <= WPIPE_ConvTranspose_output_pipe_580_inst_req_1;
      update_req_unguarded(45) <= WPIPE_ConvTranspose_output_pipe_774_inst_req_1;
      update_req_unguarded(44) <= WPIPE_ConvTranspose_output_pipe_543_inst_req_1;
      update_req_unguarded(43) <= WPIPE_ConvTranspose_output_pipe_601_inst_req_1;
      update_req_unguarded(42) <= WPIPE_ConvTranspose_output_pipe_685_inst_req_1;
      update_req_unguarded(41) <= WPIPE_ConvTranspose_output_pipe_622_inst_req_1;
      update_req_unguarded(40) <= WPIPE_ConvTranspose_output_pipe_37_inst_req_1;
      update_req_unguarded(39) <= WPIPE_ConvTranspose_output_pipe_643_inst_req_1;
      update_req_unguarded(38) <= WPIPE_ConvTranspose_output_pipe_664_inst_req_1;
      update_req_unguarded(37) <= WPIPE_ConvTranspose_output_pipe_874_inst_req_1;
      update_req_unguarded(36) <= WPIPE_ConvTranspose_output_pipe_811_inst_req_1;
      update_req_unguarded(35) <= WPIPE_ConvTranspose_output_pipe_559_inst_req_1;
      update_req_unguarded(34) <= WPIPE_ConvTranspose_output_pipe_832_inst_req_1;
      update_req_unguarded(33) <= WPIPE_ConvTranspose_output_pipe_853_inst_req_1;
      update_req_unguarded(32) <= WPIPE_ConvTranspose_output_pipe_895_inst_req_1;
      update_req_unguarded(31) <= WPIPE_ConvTranspose_output_pipe_916_inst_req_1;
      update_req_unguarded(30) <= WPIPE_ConvTranspose_output_pipe_53_inst_req_1;
      update_req_unguarded(29) <= WPIPE_ConvTranspose_output_pipe_68_inst_req_1;
      update_req_unguarded(28) <= WPIPE_ConvTranspose_output_pipe_84_inst_req_1;
      update_req_unguarded(27) <= WPIPE_ConvTranspose_output_pipe_99_inst_req_1;
      update_req_unguarded(26) <= WPIPE_ConvTranspose_output_pipe_115_inst_req_1;
      update_req_unguarded(25) <= WPIPE_ConvTranspose_output_pipe_130_inst_req_1;
      update_req_unguarded(24) <= WPIPE_ConvTranspose_output_pipe_146_inst_req_1;
      update_req_unguarded(23) <= WPIPE_ConvTranspose_output_pipe_161_inst_req_1;
      update_req_unguarded(22) <= WPIPE_ConvTranspose_output_pipe_177_inst_req_1;
      update_req_unguarded(21) <= WPIPE_ConvTranspose_output_pipe_192_inst_req_1;
      update_req_unguarded(20) <= WPIPE_ConvTranspose_output_pipe_208_inst_req_1;
      update_req_unguarded(19) <= WPIPE_ConvTranspose_output_pipe_223_inst_req_1;
      update_req_unguarded(18) <= WPIPE_ConvTranspose_output_pipe_239_inst_req_1;
      update_req_unguarded(17) <= WPIPE_ConvTranspose_output_pipe_307_inst_req_1;
      update_req_unguarded(16) <= WPIPE_ConvTranspose_output_pipe_323_inst_req_1;
      update_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_338_inst_req_1;
      update_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_354_inst_req_1;
      update_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_369_inst_req_1;
      update_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_385_inst_req_1;
      update_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_400_inst_req_1;
      update_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_416_inst_req_1;
      update_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_431_inst_req_1;
      update_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_447_inst_req_1;
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1383_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1386_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1389_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1392_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1395_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1398_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1401_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1404_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_790_inst_ack_1 <= update_ack_unguarded(47);
      WPIPE_ConvTranspose_output_pipe_580_inst_ack_1 <= update_ack_unguarded(46);
      WPIPE_ConvTranspose_output_pipe_774_inst_ack_1 <= update_ack_unguarded(45);
      WPIPE_ConvTranspose_output_pipe_543_inst_ack_1 <= update_ack_unguarded(44);
      WPIPE_ConvTranspose_output_pipe_601_inst_ack_1 <= update_ack_unguarded(43);
      WPIPE_ConvTranspose_output_pipe_685_inst_ack_1 <= update_ack_unguarded(42);
      WPIPE_ConvTranspose_output_pipe_622_inst_ack_1 <= update_ack_unguarded(41);
      WPIPE_ConvTranspose_output_pipe_37_inst_ack_1 <= update_ack_unguarded(40);
      WPIPE_ConvTranspose_output_pipe_643_inst_ack_1 <= update_ack_unguarded(39);
      WPIPE_ConvTranspose_output_pipe_664_inst_ack_1 <= update_ack_unguarded(38);
      WPIPE_ConvTranspose_output_pipe_874_inst_ack_1 <= update_ack_unguarded(37);
      WPIPE_ConvTranspose_output_pipe_811_inst_ack_1 <= update_ack_unguarded(36);
      WPIPE_ConvTranspose_output_pipe_559_inst_ack_1 <= update_ack_unguarded(35);
      WPIPE_ConvTranspose_output_pipe_832_inst_ack_1 <= update_ack_unguarded(34);
      WPIPE_ConvTranspose_output_pipe_853_inst_ack_1 <= update_ack_unguarded(33);
      WPIPE_ConvTranspose_output_pipe_895_inst_ack_1 <= update_ack_unguarded(32);
      WPIPE_ConvTranspose_output_pipe_916_inst_ack_1 <= update_ack_unguarded(31);
      WPIPE_ConvTranspose_output_pipe_53_inst_ack_1 <= update_ack_unguarded(30);
      WPIPE_ConvTranspose_output_pipe_68_inst_ack_1 <= update_ack_unguarded(29);
      WPIPE_ConvTranspose_output_pipe_84_inst_ack_1 <= update_ack_unguarded(28);
      WPIPE_ConvTranspose_output_pipe_99_inst_ack_1 <= update_ack_unguarded(27);
      WPIPE_ConvTranspose_output_pipe_115_inst_ack_1 <= update_ack_unguarded(26);
      WPIPE_ConvTranspose_output_pipe_130_inst_ack_1 <= update_ack_unguarded(25);
      WPIPE_ConvTranspose_output_pipe_146_inst_ack_1 <= update_ack_unguarded(24);
      WPIPE_ConvTranspose_output_pipe_161_inst_ack_1 <= update_ack_unguarded(23);
      WPIPE_ConvTranspose_output_pipe_177_inst_ack_1 <= update_ack_unguarded(22);
      WPIPE_ConvTranspose_output_pipe_192_inst_ack_1 <= update_ack_unguarded(21);
      WPIPE_ConvTranspose_output_pipe_208_inst_ack_1 <= update_ack_unguarded(20);
      WPIPE_ConvTranspose_output_pipe_223_inst_ack_1 <= update_ack_unguarded(19);
      WPIPE_ConvTranspose_output_pipe_239_inst_ack_1 <= update_ack_unguarded(18);
      WPIPE_ConvTranspose_output_pipe_307_inst_ack_1 <= update_ack_unguarded(17);
      WPIPE_ConvTranspose_output_pipe_323_inst_ack_1 <= update_ack_unguarded(16);
      WPIPE_ConvTranspose_output_pipe_338_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_354_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_369_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_385_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_400_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_416_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_431_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_447_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1383_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1386_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1389_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1392_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1395_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1398_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1401_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1404_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      guard_vector(40)  <=  '1';
      guard_vector(41)  <=  '1';
      guard_vector(42)  <=  '1';
      guard_vector(43)  <=  '1';
      guard_vector(44)  <=  '1';
      guard_vector(45)  <=  '1';
      guard_vector(46)  <=  '1';
      guard_vector(47)  <=  '1';
      data_in <= call321_789 & call243_579 & call313_773 & call225_542 & call253_600 & call293_684 & call263_621 & call_36 & call273_642 & call283_663 & call361_873 & call331_810 & call233_558 & call341_831 & call351_852 & call371_894 & call381_915 & call6_52 & call13_67 & call22_83 & call30_98 & call39_114 & call47_129 & call56_145 & call64_160 & call73_176 & call81_191 & call90_207 & call98_222 & call107_238 & call135_306 & call144_322 & call152_337 & call161_353 & call169_368 & call178_384 & call186_399 & call195_415 & call203_430 & call212_446 & conv541_1382 & conv535_1372 & conv529_1362 & conv523_1352 & conv517_1342 & conv511_1332 & conv505_1322 & conv499_1312;
      ConvTranspose_output_pipe_write_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_4_gI", nreqs => 48, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_4: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 48, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared outport operator group (5) : WPIPE_elapsed_time_pipe_1242_inst 
    OutportGroup_5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1242_inst_req_0;
      WPIPE_elapsed_time_pipe_1242_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1242_inst_req_1;
      WPIPE_elapsed_time_pipe_1242_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub_1241;
      elapsed_time_pipe_write_5_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_5: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 5
    -- shared call operator group (0) : call_stmt_1066_call call_stmt_1231_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1066_call_req_0;
      reqL_unguarded(0) <= call_stmt_1231_call_req_0;
      call_stmt_1066_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1231_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1066_call_req_1;
      reqR_unguarded(0) <= call_stmt_1231_call_req_1;
      call_stmt_1066_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1231_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call419_1066 <= data_out(127 downto 64);
      call478_1231 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_3912_start: Boolean;
  signal convTransposeA_CP_3912_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block0_start_1452_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1437_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1437_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1455_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1452_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1443_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1437_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1434_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1458_inst_ack_1 : boolean;
  signal type_cast_1531_inst_ack_0 : boolean;
  signal type_cast_1531_inst_req_1 : boolean;
  signal type_cast_1531_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1467_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1443_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1440_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1440_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1434_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1452_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1455_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1452_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1437_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1440_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1464_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1440_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1467_inst_ack_1 : boolean;
  signal type_cast_1591_inst_req_0 : boolean;
  signal type_cast_1591_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1464_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1467_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1467_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1449_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1461_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1434_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1443_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1449_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1461_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1458_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1464_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1434_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1449_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1464_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1443_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1458_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1449_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1461_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1446_inst_req_0 : boolean;
  signal phi_stmt_1525_ack_0 : boolean;
  signal RPIPE_Block0_start_1446_inst_ack_0 : boolean;
  signal type_cast_1591_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1446_inst_req_1 : boolean;
  signal type_cast_1591_inst_ack_0 : boolean;
  signal phi_stmt_1585_req_1 : boolean;
  signal RPIPE_Block0_start_1455_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1446_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1455_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1461_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1458_inst_req_1 : boolean;
  signal phi_stmt_1585_req_0 : boolean;
  signal type_cast_1531_inst_ack_1 : boolean;
  signal phi_stmt_1525_req_1 : boolean;
  signal phi_stmt_1585_ack_0 : boolean;
  signal type_cast_1472_inst_req_0 : boolean;
  signal type_cast_1472_inst_ack_0 : boolean;
  signal phi_stmt_1518_ack_0 : boolean;
  signal type_cast_1472_inst_req_1 : boolean;
  signal type_cast_1472_inst_ack_1 : boolean;
  signal type_cast_1476_inst_req_0 : boolean;
  signal type_cast_1476_inst_ack_0 : boolean;
  signal type_cast_1476_inst_req_1 : boolean;
  signal type_cast_1476_inst_ack_1 : boolean;
  signal type_cast_1486_inst_req_0 : boolean;
  signal type_cast_1486_inst_ack_0 : boolean;
  signal type_cast_1486_inst_req_1 : boolean;
  signal type_cast_1486_inst_ack_1 : boolean;
  signal type_cast_1613_inst_req_0 : boolean;
  signal type_cast_1613_inst_ack_0 : boolean;
  signal type_cast_1613_inst_req_1 : boolean;
  signal type_cast_1613_inst_ack_1 : boolean;
  signal type_cast_1627_inst_req_0 : boolean;
  signal type_cast_1627_inst_ack_0 : boolean;
  signal type_cast_1627_inst_req_1 : boolean;
  signal type_cast_1627_inst_ack_1 : boolean;
  signal array_obj_ref_1633_index_offset_req_0 : boolean;
  signal array_obj_ref_1633_index_offset_ack_0 : boolean;
  signal array_obj_ref_1633_index_offset_req_1 : boolean;
  signal array_obj_ref_1633_index_offset_ack_1 : boolean;
  signal addr_of_1634_final_reg_req_0 : boolean;
  signal addr_of_1634_final_reg_ack_0 : boolean;
  signal addr_of_1634_final_reg_req_1 : boolean;
  signal addr_of_1634_final_reg_ack_1 : boolean;
  signal ptr_deref_1638_load_0_req_0 : boolean;
  signal ptr_deref_1638_load_0_ack_0 : boolean;
  signal ptr_deref_1638_load_0_req_1 : boolean;
  signal ptr_deref_1638_load_0_ack_1 : boolean;
  signal type_cast_1643_inst_req_0 : boolean;
  signal type_cast_1643_inst_ack_0 : boolean;
  signal type_cast_1643_inst_req_1 : boolean;
  signal type_cast_1643_inst_ack_1 : boolean;
  signal type_cast_1657_inst_req_0 : boolean;
  signal type_cast_1657_inst_ack_0 : boolean;
  signal type_cast_1657_inst_req_1 : boolean;
  signal type_cast_1657_inst_ack_1 : boolean;
  signal array_obj_ref_1663_index_offset_req_0 : boolean;
  signal array_obj_ref_1663_index_offset_ack_0 : boolean;
  signal array_obj_ref_1663_index_offset_req_1 : boolean;
  signal array_obj_ref_1663_index_offset_ack_1 : boolean;
  signal addr_of_1664_final_reg_req_0 : boolean;
  signal addr_of_1664_final_reg_ack_0 : boolean;
  signal addr_of_1664_final_reg_req_1 : boolean;
  signal addr_of_1664_final_reg_ack_1 : boolean;
  signal ptr_deref_1667_store_0_req_0 : boolean;
  signal ptr_deref_1667_store_0_ack_0 : boolean;
  signal ptr_deref_1667_store_0_req_1 : boolean;
  signal ptr_deref_1667_store_0_ack_1 : boolean;
  signal type_cast_1673_inst_req_0 : boolean;
  signal type_cast_1673_inst_ack_0 : boolean;
  signal type_cast_1673_inst_req_1 : boolean;
  signal type_cast_1673_inst_ack_1 : boolean;
  signal if_stmt_1688_branch_req_0 : boolean;
  signal if_stmt_1688_branch_ack_1 : boolean;
  signal if_stmt_1688_branch_ack_0 : boolean;
  signal type_cast_1712_inst_req_0 : boolean;
  signal type_cast_1712_inst_ack_0 : boolean;
  signal type_cast_1712_inst_req_1 : boolean;
  signal type_cast_1712_inst_ack_1 : boolean;
  signal type_cast_1721_inst_req_0 : boolean;
  signal type_cast_1721_inst_ack_0 : boolean;
  signal type_cast_1721_inst_req_1 : boolean;
  signal type_cast_1721_inst_ack_1 : boolean;
  signal type_cast_1738_inst_req_0 : boolean;
  signal type_cast_1738_inst_ack_0 : boolean;
  signal type_cast_1738_inst_req_1 : boolean;
  signal type_cast_1738_inst_ack_1 : boolean;
  signal if_stmt_1745_branch_req_0 : boolean;
  signal if_stmt_1745_branch_ack_1 : boolean;
  signal if_stmt_1745_branch_ack_0 : boolean;
  signal WPIPE_Block0_done_1753_inst_req_0 : boolean;
  signal WPIPE_Block0_done_1753_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1753_inst_req_1 : boolean;
  signal WPIPE_Block0_done_1753_inst_ack_1 : boolean;
  signal phi_stmt_1518_req_0 : boolean;
  signal phi_stmt_1525_req_0 : boolean;
  signal type_cast_1524_inst_req_0 : boolean;
  signal type_cast_1524_inst_ack_0 : boolean;
  signal type_cast_1524_inst_req_1 : boolean;
  signal type_cast_1524_inst_ack_1 : boolean;
  signal phi_stmt_1518_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_3912_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3912_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_3912_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3912_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_3912: Block -- control-path 
    signal convTransposeA_CP_3912_elements: BooleanArray(87 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_3912_elements(0) <= convTransposeA_CP_3912_start;
    convTransposeA_CP_3912_symbol <= convTransposeA_CP_3912_elements(67);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_1432/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1434_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468__entry__
      -- CP-element group 0: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1434_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1432/branch_block_stmt_1432__entry__
      -- CP-element group 0: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1434_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/$entry
      -- 
    rr_3960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(0), ack => RPIPE_Block0_start_1434_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1434_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1434_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1434_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1434_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1434_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1434_Update/cr
      -- 
    ra_3961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1434_inst_ack_0, ack => convTransposeA_CP_3912_elements(1)); -- 
    cr_3965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(1), ack => RPIPE_Block0_start_1434_inst_req_1); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1437_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1434_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1434_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1434_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1437_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1437_Sample/$entry
      -- 
    ca_3966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1434_inst_ack_1, ack => convTransposeA_CP_3912_elements(2)); -- 
    rr_3974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(2), ack => RPIPE_Block0_start_1437_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1437_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1437_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1437_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1437_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1437_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1437_update_start_
      -- 
    ra_3975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1437_inst_ack_0, ack => convTransposeA_CP_3912_elements(3)); -- 
    cr_3979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(3), ack => RPIPE_Block0_start_1437_inst_req_1); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1437_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1440_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1440_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1440_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1437_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1437_update_completed_
      -- 
    ca_3980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1437_inst_ack_1, ack => convTransposeA_CP_3912_elements(4)); -- 
    rr_3988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(4), ack => RPIPE_Block0_start_1440_inst_req_0); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1440_update_start_
      -- CP-element group 5: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1440_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1440_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1440_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1440_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1440_Update/cr
      -- 
    ra_3989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1440_inst_ack_0, ack => convTransposeA_CP_3912_elements(5)); -- 
    cr_3993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(5), ack => RPIPE_Block0_start_1440_inst_req_1); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1440_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1440_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1440_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1443_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1443_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1443_Sample/rr
      -- 
    ca_3994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1440_inst_ack_1, ack => convTransposeA_CP_3912_elements(6)); -- 
    rr_4002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(6), ack => RPIPE_Block0_start_1443_inst_req_0); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1443_Update/cr
      -- CP-element group 7: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1443_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1443_update_start_
      -- CP-element group 7: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1443_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1443_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1443_Update/$entry
      -- 
    ra_4003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1443_inst_ack_0, ack => convTransposeA_CP_3912_elements(7)); -- 
    cr_4007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(7), ack => RPIPE_Block0_start_1443_inst_req_1); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1443_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1446_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1443_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1446_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1446_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1443_Update/$exit
      -- 
    ca_4008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1443_inst_ack_1, ack => convTransposeA_CP_3912_elements(8)); -- 
    rr_4016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(8), ack => RPIPE_Block0_start_1446_inst_req_0); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1446_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1446_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1446_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1446_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1446_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1446_Update/cr
      -- 
    ra_4017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1446_inst_ack_0, ack => convTransposeA_CP_3912_elements(9)); -- 
    cr_4021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(9), ack => RPIPE_Block0_start_1446_inst_req_1); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1449_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1449_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1446_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1446_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1446_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1449_sample_start_
      -- 
    ca_4022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1446_inst_ack_1, ack => convTransposeA_CP_3912_elements(10)); -- 
    rr_4030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(10), ack => RPIPE_Block0_start_1449_inst_req_0); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1449_update_start_
      -- CP-element group 11: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1449_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1449_Update/cr
      -- CP-element group 11: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1449_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1449_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1449_sample_completed_
      -- 
    ra_4031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1449_inst_ack_0, ack => convTransposeA_CP_3912_elements(11)); -- 
    cr_4035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(11), ack => RPIPE_Block0_start_1449_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1449_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1452_Sample/rr
      -- CP-element group 12: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1452_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1449_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1449_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1452_Sample/$entry
      -- 
    ca_4036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1449_inst_ack_1, ack => convTransposeA_CP_3912_elements(12)); -- 
    rr_4044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(12), ack => RPIPE_Block0_start_1452_inst_req_0); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1452_Update/cr
      -- CP-element group 13: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1452_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1452_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1452_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1452_update_start_
      -- CP-element group 13: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1452_Sample/$exit
      -- 
    ra_4045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1452_inst_ack_0, ack => convTransposeA_CP_3912_elements(13)); -- 
    cr_4049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(13), ack => RPIPE_Block0_start_1452_inst_req_1); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1452_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1452_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1455_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1452_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1455_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1455_Sample/rr
      -- 
    ca_4050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1452_inst_ack_1, ack => convTransposeA_CP_3912_elements(14)); -- 
    rr_4058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(14), ack => RPIPE_Block0_start_1455_inst_req_0); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1455_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1455_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1455_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1455_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1455_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1455_Sample/ra
      -- 
    ra_4059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1455_inst_ack_0, ack => convTransposeA_CP_3912_elements(15)); -- 
    cr_4063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(15), ack => RPIPE_Block0_start_1455_inst_req_1); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1455_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1458_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1458_Sample/rr
      -- CP-element group 16: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1455_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1455_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1458_sample_start_
      -- 
    ca_4064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1455_inst_ack_1, ack => convTransposeA_CP_3912_elements(16)); -- 
    rr_4072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(16), ack => RPIPE_Block0_start_1458_inst_req_0); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1458_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1458_update_start_
      -- CP-element group 17: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1458_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1458_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1458_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1458_Update/cr
      -- 
    ra_4073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1458_inst_ack_0, ack => convTransposeA_CP_3912_elements(17)); -- 
    cr_4077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(17), ack => RPIPE_Block0_start_1458_inst_req_1); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1458_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1458_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1461_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1461_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1461_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1458_Update/$exit
      -- 
    ca_4078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1458_inst_ack_1, ack => convTransposeA_CP_3912_elements(18)); -- 
    rr_4086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(18), ack => RPIPE_Block0_start_1461_inst_req_0); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1461_Update/cr
      -- CP-element group 19: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1461_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1461_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1461_update_start_
      -- CP-element group 19: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1461_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1461_Sample/$exit
      -- 
    ra_4087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1461_inst_ack_0, ack => convTransposeA_CP_3912_elements(19)); -- 
    cr_4091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(19), ack => RPIPE_Block0_start_1461_inst_req_1); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1464_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1461_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1464_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1461_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1461_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1464_sample_start_
      -- 
    ca_4092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1461_inst_ack_1, ack => convTransposeA_CP_3912_elements(20)); -- 
    rr_4100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(20), ack => RPIPE_Block0_start_1464_inst_req_0); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1464_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1464_Update/cr
      -- CP-element group 21: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1464_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1464_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1464_update_start_
      -- CP-element group 21: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1464_Update/$entry
      -- 
    ra_4101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1464_inst_ack_0, ack => convTransposeA_CP_3912_elements(21)); -- 
    cr_4105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(21), ack => RPIPE_Block0_start_1464_inst_req_1); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1467_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1467_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1467_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1464_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1464_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1464_Update/$exit
      -- 
    ca_4106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1464_inst_ack_1, ack => convTransposeA_CP_3912_elements(22)); -- 
    rr_4114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(22), ack => RPIPE_Block0_start_1467_inst_req_0); -- 
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1467_Update/cr
      -- CP-element group 23: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1467_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1467_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1467_update_start_
      -- CP-element group 23: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1467_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1467_Sample/ra
      -- 
    ra_4115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1467_inst_ack_0, ack => convTransposeA_CP_3912_elements(23)); -- 
    cr_4119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(23), ack => RPIPE_Block0_start_1467_inst_req_1); -- 
    -- CP-element group 24:  fork  transition  place  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	27 
    -- CP-element group 24: 	28 
    -- CP-element group 24: 	29 
    -- CP-element group 24: 	30 
    -- CP-element group 24:  members (25) 
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1467_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/$exit
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468__exit__
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515__entry__
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1467_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1435_to_assign_stmt_1468/RPIPE_Block0_start_1467_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/$entry
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1472_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1472_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1472_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1472_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1472_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1472_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1476_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1476_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1476_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1476_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1476_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1476_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1486_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1486_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1486_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1486_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1486_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1486_Update/cr
      -- 
    ca_4120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1467_inst_ack_1, ack => convTransposeA_CP_3912_elements(24)); -- 
    rr_4131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(24), ack => type_cast_1472_inst_req_0); -- 
    cr_4136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(24), ack => type_cast_1472_inst_req_1); -- 
    rr_4145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(24), ack => type_cast_1476_inst_req_0); -- 
    cr_4150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(24), ack => type_cast_1476_inst_req_1); -- 
    rr_4159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(24), ack => type_cast_1486_inst_req_0); -- 
    cr_4164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(24), ack => type_cast_1486_inst_req_1); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1472_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1472_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1472_Sample/ra
      -- 
    ra_4132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1472_inst_ack_0, ack => convTransposeA_CP_3912_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1472_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1472_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1472_Update/ca
      -- 
    ca_4137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1472_inst_ack_1, ack => convTransposeA_CP_3912_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	24 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1476_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1476_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1476_Sample/ra
      -- 
    ra_4146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1476_inst_ack_0, ack => convTransposeA_CP_3912_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	24 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1476_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1476_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1476_Update/ca
      -- 
    ca_4151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1476_inst_ack_1, ack => convTransposeA_CP_3912_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	24 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1486_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1486_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1486_Sample/ra
      -- 
    ra_4160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1486_inst_ack_0, ack => convTransposeA_CP_3912_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	24 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1486_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1486_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/type_cast_1486_Update/ca
      -- 
    ca_4165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1486_inst_ack_1, ack => convTransposeA_CP_3912_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	68 
    -- CP-element group 31: 	69 
    -- CP-element group 31:  members (8) 
      -- CP-element group 31: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515__exit__
      -- CP-element group 31: 	 branch_block_stmt_1432/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_1432/assign_stmt_1473_to_assign_stmt_1515/$exit
      -- CP-element group 31: 	 branch_block_stmt_1432/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_1432/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/$entry
      -- CP-element group 31: 	 branch_block_stmt_1432/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/phi_stmt_1518_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1432/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/$entry
      -- CP-element group 31: 	 branch_block_stmt_1432/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/phi_stmt_1525_sources/$entry
      -- 
    convTransposeA_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3912_elements(26) & convTransposeA_CP_3912_elements(28) & convTransposeA_CP_3912_elements(30);
      gj_convTransposeA_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3912_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	87 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1613_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1613_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1613_Sample/ra
      -- 
    ra_4180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1613_inst_ack_0, ack => convTransposeA_CP_3912_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	87 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1613_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1613_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1613_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1627_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1627_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1627_Sample/rr
      -- 
    ca_4185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1613_inst_ack_1, ack => convTransposeA_CP_3912_elements(33)); -- 
    rr_4193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(33), ack => type_cast_1627_inst_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1627_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1627_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1627_Sample/ra
      -- 
    ra_4194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1627_inst_ack_0, ack => convTransposeA_CP_3912_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	87 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (16) 
      -- CP-element group 35: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1627_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1627_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1627_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_index_resized_1
      -- CP-element group 35: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_index_scaled_1
      -- CP-element group 35: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_index_computed_1
      -- CP-element group 35: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_index_resize_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_index_resize_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_index_resize_1/index_resize_req
      -- CP-element group 35: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_index_resize_1/index_resize_ack
      -- CP-element group 35: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_index_scale_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_index_scale_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_index_scale_1/scale_rename_req
      -- CP-element group 35: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_index_scale_1/scale_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_final_index_sum_regn_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_final_index_sum_regn_Sample/req
      -- 
    ca_4199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1627_inst_ack_1, ack => convTransposeA_CP_3912_elements(35)); -- 
    req_4224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(35), ack => array_obj_ref_1633_index_offset_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	55 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_final_index_sum_regn_sample_complete
      -- CP-element group 36: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_final_index_sum_regn_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_final_index_sum_regn_Sample/ack
      -- 
    ack_4225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1633_index_offset_ack_0, ack => convTransposeA_CP_3912_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	87 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (11) 
      -- CP-element group 37: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1634_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_offset_calculated
      -- CP-element group 37: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_final_index_sum_regn_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_final_index_sum_regn_Update/ack
      -- CP-element group 37: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_base_plus_offset/$entry
      -- CP-element group 37: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_base_plus_offset/$exit
      -- CP-element group 37: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_base_plus_offset/sum_rename_req
      -- CP-element group 37: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1634_request/$entry
      -- CP-element group 37: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1634_request/req
      -- 
    ack_4230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1633_index_offset_ack_1, ack => convTransposeA_CP_3912_elements(37)); -- 
    req_4239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(37), ack => addr_of_1634_final_reg_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1634_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1634_request/$exit
      -- CP-element group 38: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1634_request/ack
      -- 
    ack_4240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1634_final_reg_ack_0, ack => convTransposeA_CP_3912_elements(38)); -- 
    -- CP-element group 39:  join  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	87 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (24) 
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1634_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1634_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1634_complete/ack
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_base_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_word_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_base_address_resized
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_base_addr_resize/$entry
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_base_addr_resize/$exit
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_base_addr_resize/base_resize_req
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_base_addr_resize/base_resize_ack
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_word_addrgen/$entry
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_word_addrgen/$exit
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_word_addrgen/root_register_req
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_word_addrgen/root_register_ack
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_Sample/word_access_start/$entry
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_Sample/word_access_start/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_Sample/word_access_start/word_0/rr
      -- 
    ack_4245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1634_final_reg_ack_1, ack => convTransposeA_CP_3912_elements(39)); -- 
    rr_4278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(39), ack => ptr_deref_1638_load_0_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_Sample/word_access_start/$exit
      -- CP-element group 40: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_Sample/word_access_start/word_0/$exit
      -- CP-element group 40: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_Sample/word_access_start/word_0/ra
      -- 
    ra_4279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1638_load_0_ack_0, ack => convTransposeA_CP_3912_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	87 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	50 
    -- CP-element group 41:  members (9) 
      -- CP-element group 41: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_Update/word_access_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_Update/word_access_complete/word_0/$exit
      -- CP-element group 41: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_Update/word_access_complete/word_0/ca
      -- CP-element group 41: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_Update/ptr_deref_1638_Merge/$entry
      -- CP-element group 41: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_Update/ptr_deref_1638_Merge/$exit
      -- CP-element group 41: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_Update/ptr_deref_1638_Merge/merge_req
      -- CP-element group 41: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_Update/ptr_deref_1638_Merge/merge_ack
      -- 
    ca_4290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1638_load_0_ack_1, ack => convTransposeA_CP_3912_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	87 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1643_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1643_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1643_Sample/ra
      -- 
    ra_4304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1643_inst_ack_0, ack => convTransposeA_CP_3912_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	87 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1643_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1643_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1643_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1657_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1657_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1657_Sample/rr
      -- 
    ca_4309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1643_inst_ack_1, ack => convTransposeA_CP_3912_elements(43)); -- 
    rr_4317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(43), ack => type_cast_1657_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1657_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1657_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1657_Sample/ra
      -- 
    ra_4318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1657_inst_ack_0, ack => convTransposeA_CP_3912_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	87 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (16) 
      -- CP-element group 45: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1657_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1657_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1657_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_index_resized_1
      -- CP-element group 45: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_index_scaled_1
      -- CP-element group 45: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_index_computed_1
      -- CP-element group 45: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_index_resize_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_index_resize_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_index_resize_1/index_resize_req
      -- CP-element group 45: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_index_resize_1/index_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_index_scale_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_index_scale_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_index_scale_1/scale_rename_req
      -- CP-element group 45: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_index_scale_1/scale_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_final_index_sum_regn_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_final_index_sum_regn_Sample/req
      -- 
    ca_4323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1657_inst_ack_1, ack => convTransposeA_CP_3912_elements(45)); -- 
    req_4348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(45), ack => array_obj_ref_1663_index_offset_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	55 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_final_index_sum_regn_sample_complete
      -- CP-element group 46: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_final_index_sum_regn_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_final_index_sum_regn_Sample/ack
      -- 
    ack_4349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1663_index_offset_ack_0, ack => convTransposeA_CP_3912_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	87 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (11) 
      -- CP-element group 47: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1664_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_root_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_offset_calculated
      -- CP-element group 47: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_final_index_sum_regn_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_final_index_sum_regn_Update/ack
      -- CP-element group 47: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_base_plus_offset/$entry
      -- CP-element group 47: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_base_plus_offset/$exit
      -- CP-element group 47: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_base_plus_offset/sum_rename_req
      -- CP-element group 47: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_base_plus_offset/sum_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1664_request/$entry
      -- CP-element group 47: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1664_request/req
      -- 
    ack_4354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1663_index_offset_ack_1, ack => convTransposeA_CP_3912_elements(47)); -- 
    req_4363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(47), ack => addr_of_1664_final_reg_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1664_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1664_request/$exit
      -- CP-element group 48: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1664_request/ack
      -- 
    ack_4364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1664_final_reg_ack_0, ack => convTransposeA_CP_3912_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	87 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (19) 
      -- CP-element group 49: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1664_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1664_complete/$exit
      -- CP-element group 49: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1664_complete/ack
      -- CP-element group 49: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_base_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_word_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_base_address_resized
      -- CP-element group 49: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_base_addr_resize/$entry
      -- CP-element group 49: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_base_addr_resize/$exit
      -- CP-element group 49: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_base_addr_resize/base_resize_req
      -- CP-element group 49: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_base_addr_resize/base_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_word_addrgen/$entry
      -- CP-element group 49: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_word_addrgen/$exit
      -- CP-element group 49: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_word_addrgen/root_register_req
      -- CP-element group 49: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_word_addrgen/root_register_ack
      -- 
    ack_4369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1664_final_reg_ack_1, ack => convTransposeA_CP_3912_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: 	41 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_Sample/ptr_deref_1667_Split/$entry
      -- CP-element group 50: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_Sample/ptr_deref_1667_Split/$exit
      -- CP-element group 50: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_Sample/ptr_deref_1667_Split/split_req
      -- CP-element group 50: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_Sample/ptr_deref_1667_Split/split_ack
      -- CP-element group 50: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_Sample/word_access_start/$entry
      -- CP-element group 50: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_Sample/word_access_start/word_0/$entry
      -- CP-element group 50: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_Sample/word_access_start/word_0/rr
      -- 
    rr_4407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(50), ack => ptr_deref_1667_store_0_req_0); -- 
    convTransposeA_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3912_elements(49) & convTransposeA_CP_3912_elements(41);
      gj_convTransposeA_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3912_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_Sample/word_access_start/$exit
      -- CP-element group 51: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_Sample/word_access_start/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_Sample/word_access_start/word_0/ra
      -- 
    ra_4408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1667_store_0_ack_0, ack => convTransposeA_CP_3912_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	87 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_Update/word_access_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_Update/word_access_complete/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_Update/word_access_complete/word_0/ca
      -- 
    ca_4419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1667_store_0_ack_1, ack => convTransposeA_CP_3912_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	87 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1673_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1673_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1673_Sample/ra
      -- 
    ra_4428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1673_inst_ack_0, ack => convTransposeA_CP_3912_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	87 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1673_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1673_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1673_Update/ca
      -- 
    ca_4433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1673_inst_ack_1, ack => convTransposeA_CP_3912_elements(54)); -- 
    -- CP-element group 55:  branch  join  transition  place  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	36 
    -- CP-element group 55: 	46 
    -- CP-element group 55: 	54 
    -- CP-element group 55: 	52 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (10) 
      -- CP-element group 55: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687__exit__
      -- CP-element group 55: 	 branch_block_stmt_1432/if_stmt_1688__entry__
      -- CP-element group 55: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/$exit
      -- CP-element group 55: 	 branch_block_stmt_1432/if_stmt_1688_dead_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_1432/if_stmt_1688_eval_test/$entry
      -- CP-element group 55: 	 branch_block_stmt_1432/if_stmt_1688_eval_test/$exit
      -- CP-element group 55: 	 branch_block_stmt_1432/if_stmt_1688_eval_test/branch_req
      -- CP-element group 55: 	 branch_block_stmt_1432/R_cmp_1689_place
      -- CP-element group 55: 	 branch_block_stmt_1432/if_stmt_1688_if_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_1432/if_stmt_1688_else_link/$entry
      -- 
    branch_req_4441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(55), ack => if_stmt_1688_branch_req_0); -- 
    convTransposeA_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3912_elements(36) & convTransposeA_CP_3912_elements(46) & convTransposeA_CP_3912_elements(54) & convTransposeA_CP_3912_elements(52);
      gj_convTransposeA_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3912_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	82 
    -- CP-element group 56: 	83 
    -- CP-element group 56:  members (24) 
      -- CP-element group 56: 	 branch_block_stmt_1432/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_1432/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_1432/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1585/$entry
      -- CP-element group 56: 	 branch_block_stmt_1432/merge_stmt_1694_PhiAck/$exit
      -- CP-element group 56: 	 branch_block_stmt_1432/merge_stmt_1694_PhiAck/$entry
      -- CP-element group 56: 	 branch_block_stmt_1432/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_1432/merge_stmt_1694_PhiReqMerge
      -- CP-element group 56: 	 branch_block_stmt_1432/merge_stmt_1694__exit__
      -- CP-element group 56: 	 branch_block_stmt_1432/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1585/phi_stmt_1585_sources/type_cast_1591/SplitProtocol/Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_1432/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1585/phi_stmt_1585_sources/type_cast_1591/SplitProtocol/Update/cr
      -- CP-element group 56: 	 branch_block_stmt_1432/assign_stmt_1700__entry__
      -- CP-element group 56: 	 branch_block_stmt_1432/assign_stmt_1700__exit__
      -- CP-element group 56: 	 branch_block_stmt_1432/ifx_xthen_whilex_xbody
      -- CP-element group 56: 	 branch_block_stmt_1432/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1585/phi_stmt_1585_sources/type_cast_1591/SplitProtocol/Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_1432/merge_stmt_1694_PhiAck/dummy
      -- CP-element group 56: 	 branch_block_stmt_1432/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1585/phi_stmt_1585_sources/$entry
      -- CP-element group 56: 	 branch_block_stmt_1432/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1585/phi_stmt_1585_sources/type_cast_1591/SplitProtocol/Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_1432/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1585/phi_stmt_1585_sources/type_cast_1591/SplitProtocol/$entry
      -- CP-element group 56: 	 branch_block_stmt_1432/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1585/phi_stmt_1585_sources/type_cast_1591/$entry
      -- CP-element group 56: 	 branch_block_stmt_1432/if_stmt_1688_if_link/$exit
      -- CP-element group 56: 	 branch_block_stmt_1432/if_stmt_1688_if_link/if_choice_transition
      -- CP-element group 56: 	 branch_block_stmt_1432/whilex_xbody_ifx_xthen
      -- CP-element group 56: 	 branch_block_stmt_1432/assign_stmt_1700/$entry
      -- CP-element group 56: 	 branch_block_stmt_1432/assign_stmt_1700/$exit
      -- 
    if_choice_transition_4446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1688_branch_ack_1, ack => convTransposeA_CP_3912_elements(56)); -- 
    rr_4629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(56), ack => type_cast_1591_inst_req_0); -- 
    cr_4634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(56), ack => type_cast_1591_inst_req_1); -- 
    -- CP-element group 57:  fork  transition  place  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	59 
    -- CP-element group 57: 	61 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (24) 
      -- CP-element group 57: 	 branch_block_stmt_1432/merge_stmt_1702_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_1432/merge_stmt_1702__exit__
      -- CP-element group 57: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744__entry__
      -- CP-element group 57: 	 branch_block_stmt_1432/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_1432/merge_stmt_1702_PhiAck/dummy
      -- CP-element group 57: 	 branch_block_stmt_1432/merge_stmt_1702_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_1432/merge_stmt_1702_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_1432/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_1432/if_stmt_1688_else_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_1432/if_stmt_1688_else_link/else_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_1432/whilex_xbody_ifx_xelse
      -- CP-element group 57: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/$entry
      -- CP-element group 57: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1712_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1712_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1712_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1712_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1712_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1712_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1721_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1721_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1721_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1738_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1738_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1738_Update/cr
      -- 
    else_choice_transition_4450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1688_branch_ack_0, ack => convTransposeA_CP_3912_elements(57)); -- 
    rr_4466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(57), ack => type_cast_1712_inst_req_0); -- 
    cr_4471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(57), ack => type_cast_1712_inst_req_1); -- 
    cr_4485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(57), ack => type_cast_1721_inst_req_1); -- 
    cr_4499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(57), ack => type_cast_1738_inst_req_1); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1712_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1712_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1712_Sample/ra
      -- 
    ra_4467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1712_inst_ack_0, ack => convTransposeA_CP_3912_elements(58)); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1712_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1712_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1712_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1721_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1721_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1721_Sample/rr
      -- 
    ca_4472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1712_inst_ack_1, ack => convTransposeA_CP_3912_elements(59)); -- 
    rr_4480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(59), ack => type_cast_1721_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1721_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1721_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1721_Sample/ra
      -- 
    ra_4481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1721_inst_ack_0, ack => convTransposeA_CP_3912_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	57 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1721_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1721_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1721_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1738_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1738_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1738_Sample/rr
      -- 
    ca_4486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1721_inst_ack_1, ack => convTransposeA_CP_3912_elements(61)); -- 
    rr_4494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(61), ack => type_cast_1738_inst_req_0); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1738_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1738_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1738_Sample/ra
      -- 
    ra_4495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1738_inst_ack_0, ack => convTransposeA_CP_3912_elements(62)); -- 
    -- CP-element group 63:  branch  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (13) 
      -- CP-element group 63: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744__exit__
      -- CP-element group 63: 	 branch_block_stmt_1432/if_stmt_1745__entry__
      -- CP-element group 63: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/$exit
      -- CP-element group 63: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1738_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1738_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_1432/assign_stmt_1708_to_assign_stmt_1744/type_cast_1738_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_1432/if_stmt_1745_dead_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1432/if_stmt_1745_eval_test/$entry
      -- CP-element group 63: 	 branch_block_stmt_1432/if_stmt_1745_eval_test/$exit
      -- CP-element group 63: 	 branch_block_stmt_1432/if_stmt_1745_eval_test/branch_req
      -- CP-element group 63: 	 branch_block_stmt_1432/R_cmp116_1746_place
      -- CP-element group 63: 	 branch_block_stmt_1432/if_stmt_1745_if_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1432/if_stmt_1745_else_link/$entry
      -- 
    ca_4500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1738_inst_ack_1, ack => convTransposeA_CP_3912_elements(63)); -- 
    branch_req_4508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(63), ack => if_stmt_1745_branch_req_0); -- 
    -- CP-element group 64:  merge  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (15) 
      -- CP-element group 64: 	 branch_block_stmt_1432/merge_stmt_1751_PhiAck/dummy
      -- CP-element group 64: 	 branch_block_stmt_1432/assign_stmt_1756__entry__
      -- CP-element group 64: 	 branch_block_stmt_1432/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 64: 	 branch_block_stmt_1432/merge_stmt_1751_PhiReqMerge
      -- CP-element group 64: 	 branch_block_stmt_1432/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_1432/merge_stmt_1751_PhiAck/$entry
      -- CP-element group 64: 	 branch_block_stmt_1432/merge_stmt_1751_PhiAck/$exit
      -- CP-element group 64: 	 branch_block_stmt_1432/merge_stmt_1751__exit__
      -- CP-element group 64: 	 branch_block_stmt_1432/if_stmt_1745_if_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_1432/if_stmt_1745_if_link/if_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_1432/ifx_xelse_whilex_xend
      -- CP-element group 64: 	 branch_block_stmt_1432/assign_stmt_1756/$entry
      -- CP-element group 64: 	 branch_block_stmt_1432/assign_stmt_1756/WPIPE_Block0_done_1753_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_1432/assign_stmt_1756/WPIPE_Block0_done_1753_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1432/assign_stmt_1756/WPIPE_Block0_done_1753_Sample/req
      -- 
    if_choice_transition_4513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1745_branch_ack_1, ack => convTransposeA_CP_3912_elements(64)); -- 
    req_4530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(64), ack => WPIPE_Block0_done_1753_inst_req_0); -- 
    -- CP-element group 65:  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	71 
    -- CP-element group 65: 	72 
    -- CP-element group 65: 	74 
    -- CP-element group 65: 	75 
    -- CP-element group 65:  members (20) 
      -- CP-element group 65: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/phi_stmt_1525_sources/type_cast_1531/SplitProtocol/Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/phi_stmt_1525_sources/type_cast_1531/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/phi_stmt_1525_sources/type_cast_1531/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/phi_stmt_1525_sources/type_cast_1531/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1432/if_stmt_1745_else_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_1432/if_stmt_1745_else_link/else_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 65: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/$entry
      -- CP-element group 65: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/phi_stmt_1518_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/phi_stmt_1518_sources/type_cast_1524/$entry
      -- CP-element group 65: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/phi_stmt_1518_sources/type_cast_1524/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/phi_stmt_1518_sources/type_cast_1524/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/phi_stmt_1518_sources/type_cast_1524/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/phi_stmt_1518_sources/type_cast_1524/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/phi_stmt_1518_sources/type_cast_1524/SplitProtocol/Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/$entry
      -- CP-element group 65: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/phi_stmt_1525_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/phi_stmt_1525_sources/type_cast_1531/$entry
      -- CP-element group 65: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/phi_stmt_1525_sources/type_cast_1531/SplitProtocol/$entry
      -- 
    else_choice_transition_4517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1745_branch_ack_0, ack => convTransposeA_CP_3912_elements(65)); -- 
    cr_4602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(65), ack => type_cast_1531_inst_req_1); -- 
    rr_4597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(65), ack => type_cast_1531_inst_req_0); -- 
    rr_4574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(65), ack => type_cast_1524_inst_req_0); -- 
    cr_4579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(65), ack => type_cast_1524_inst_req_1); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_1432/assign_stmt_1756/WPIPE_Block0_done_1753_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1432/assign_stmt_1756/WPIPE_Block0_done_1753_update_start_
      -- CP-element group 66: 	 branch_block_stmt_1432/assign_stmt_1756/WPIPE_Block0_done_1753_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1432/assign_stmt_1756/WPIPE_Block0_done_1753_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_1432/assign_stmt_1756/WPIPE_Block0_done_1753_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1432/assign_stmt_1756/WPIPE_Block0_done_1753_Update/req
      -- 
    ack_4531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1753_inst_ack_0, ack => convTransposeA_CP_3912_elements(66)); -- 
    req_4535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(66), ack => WPIPE_Block0_done_1753_inst_req_1); -- 
    -- CP-element group 67:  transition  place  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (16) 
      -- CP-element group 67: 	 $exit
      -- CP-element group 67: 	 branch_block_stmt_1432/$exit
      -- CP-element group 67: 	 branch_block_stmt_1432/branch_block_stmt_1432__exit__
      -- CP-element group 67: 	 branch_block_stmt_1432/return___PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_1432/assign_stmt_1756__exit__
      -- CP-element group 67: 	 branch_block_stmt_1432/merge_stmt_1758_PhiAck/dummy
      -- CP-element group 67: 	 branch_block_stmt_1432/return__
      -- CP-element group 67: 	 branch_block_stmt_1432/merge_stmt_1758__exit__
      -- CP-element group 67: 	 branch_block_stmt_1432/merge_stmt_1758_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_1432/merge_stmt_1758_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_1432/merge_stmt_1758_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_1432/return___PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_1432/assign_stmt_1756/$exit
      -- CP-element group 67: 	 branch_block_stmt_1432/assign_stmt_1756/WPIPE_Block0_done_1753_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1432/assign_stmt_1756/WPIPE_Block0_done_1753_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1432/assign_stmt_1756/WPIPE_Block0_done_1753_Update/ack
      -- 
    ack_4536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1753_inst_ack_1, ack => convTransposeA_CP_3912_elements(67)); -- 
    -- CP-element group 68:  transition  output  delay-element  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	31 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_1432/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/$exit
      -- CP-element group 68: 	 branch_block_stmt_1432/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/phi_stmt_1518_sources/$exit
      -- CP-element group 68: 	 branch_block_stmt_1432/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/phi_stmt_1518_sources/type_cast_1522_konst_delay_trans
      -- CP-element group 68: 	 branch_block_stmt_1432/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/phi_stmt_1518_req
      -- 
    phi_stmt_1518_req_4547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1518_req_4547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(68), ack => phi_stmt_1518_req_0); -- 
    -- Element group convTransposeA_CP_3912_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => convTransposeA_CP_3912_elements(31), ack => convTransposeA_CP_3912_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  transition  output  delay-element  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	31 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_1432/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/$exit
      -- CP-element group 69: 	 branch_block_stmt_1432/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/phi_stmt_1525_sources/$exit
      -- CP-element group 69: 	 branch_block_stmt_1432/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/phi_stmt_1525_sources/type_cast_1529_konst_delay_trans
      -- CP-element group 69: 	 branch_block_stmt_1432/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/phi_stmt_1525_req
      -- 
    phi_stmt_1525_req_4555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1525_req_4555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(69), ack => phi_stmt_1525_req_0); -- 
    -- Element group convTransposeA_CP_3912_elements(69) is a control-delay.
    cp_element_69_delay: control_delay_element  generic map(name => " 69_delay", delay_value => 1)  port map(req => convTransposeA_CP_3912_elements(31), ack => convTransposeA_CP_3912_elements(69), clk => clk, reset =>reset);
    -- CP-element group 70:  join  transition  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	78 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1432/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3912_elements(68) & convTransposeA_CP_3912_elements(69);
      gj_convTransposeA_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3912_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	65 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/phi_stmt_1518_sources/type_cast_1524/SplitProtocol/Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/phi_stmt_1518_sources/type_cast_1524/SplitProtocol/Sample/ra
      -- 
    ra_4575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1524_inst_ack_0, ack => convTransposeA_CP_3912_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	65 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/phi_stmt_1518_sources/type_cast_1524/SplitProtocol/Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/phi_stmt_1518_sources/type_cast_1524/SplitProtocol/Update/ca
      -- 
    ca_4580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1524_inst_ack_1, ack => convTransposeA_CP_3912_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	77 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/$exit
      -- CP-element group 73: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/phi_stmt_1518_sources/$exit
      -- CP-element group 73: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/phi_stmt_1518_sources/type_cast_1524/$exit
      -- CP-element group 73: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/phi_stmt_1518_sources/type_cast_1524/SplitProtocol/$exit
      -- CP-element group 73: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1518/phi_stmt_1518_req
      -- 
    phi_stmt_1518_req_4581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1518_req_4581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(73), ack => phi_stmt_1518_req_1); -- 
    convTransposeA_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3912_elements(71) & convTransposeA_CP_3912_elements(72);
      gj_convTransposeA_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3912_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	65 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/phi_stmt_1525_sources/type_cast_1531/SplitProtocol/Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/phi_stmt_1525_sources/type_cast_1531/SplitProtocol/Sample/ra
      -- 
    ra_4598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1531_inst_ack_0, ack => convTransposeA_CP_3912_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	65 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/phi_stmt_1525_sources/type_cast_1531/SplitProtocol/Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/phi_stmt_1525_sources/type_cast_1531/SplitProtocol/Update/ca
      -- 
    ca_4603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1531_inst_ack_1, ack => convTransposeA_CP_3912_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/phi_stmt_1525_sources/type_cast_1531/SplitProtocol/$exit
      -- CP-element group 76: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/phi_stmt_1525_req
      -- CP-element group 76: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/$exit
      -- CP-element group 76: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/phi_stmt_1525_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1525/phi_stmt_1525_sources/type_cast_1531/$exit
      -- 
    phi_stmt_1525_req_4604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1525_req_4604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(76), ack => phi_stmt_1525_req_1); -- 
    convTransposeA_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3912_elements(74) & convTransposeA_CP_3912_elements(75);
      gj_convTransposeA_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3912_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	73 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1432/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3912_elements(73) & convTransposeA_CP_3912_elements(76);
      gj_convTransposeA_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3912_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  merge  fork  transition  place  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	70 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_1432/merge_stmt_1517_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1432/merge_stmt_1517_PhiReqMerge
      -- 
    convTransposeA_CP_3912_elements(78) <= OrReduce(convTransposeA_CP_3912_elements(70) & convTransposeA_CP_3912_elements(77));
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1432/merge_stmt_1517_PhiAck/phi_stmt_1518_ack
      -- 
    phi_stmt_1518_ack_4609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1518_ack_0, ack => convTransposeA_CP_3912_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1432/merge_stmt_1517_PhiAck/phi_stmt_1525_ack
      -- 
    phi_stmt_1525_ack_4610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1525_ack_0, ack => convTransposeA_CP_3912_elements(80)); -- 
    -- CP-element group 81:  join  transition  place  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (10) 
      -- CP-element group 81: 	 branch_block_stmt_1432/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1585/phi_stmt_1585_sources/$entry
      -- CP-element group 81: 	 branch_block_stmt_1432/merge_stmt_1517__exit__
      -- CP-element group 81: 	 branch_block_stmt_1432/assign_stmt_1537_to_assign_stmt_1582__entry__
      -- CP-element group 81: 	 branch_block_stmt_1432/assign_stmt_1537_to_assign_stmt_1582__exit__
      -- CP-element group 81: 	 branch_block_stmt_1432/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 81: 	 branch_block_stmt_1432/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1585/$entry
      -- CP-element group 81: 	 branch_block_stmt_1432/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 81: 	 branch_block_stmt_1432/merge_stmt_1517_PhiAck/$exit
      -- CP-element group 81: 	 branch_block_stmt_1432/assign_stmt_1537_to_assign_stmt_1582/$entry
      -- CP-element group 81: 	 branch_block_stmt_1432/assign_stmt_1537_to_assign_stmt_1582/$exit
      -- 
    convTransposeA_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3912_elements(79) & convTransposeA_CP_3912_elements(80);
      gj_convTransposeA_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3912_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	56 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_1432/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1585/phi_stmt_1585_sources/type_cast_1591/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_1432/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1585/phi_stmt_1585_sources/type_cast_1591/SplitProtocol/Sample/ra
      -- 
    ra_4630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1591_inst_ack_0, ack => convTransposeA_CP_3912_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	56 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1432/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1585/phi_stmt_1585_sources/type_cast_1591/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_1432/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1585/phi_stmt_1585_sources/type_cast_1591/SplitProtocol/Update/ca
      -- 
    ca_4635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1591_inst_ack_1, ack => convTransposeA_CP_3912_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (6) 
      -- CP-element group 84: 	 branch_block_stmt_1432/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 84: 	 branch_block_stmt_1432/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1585/$exit
      -- CP-element group 84: 	 branch_block_stmt_1432/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1585/phi_stmt_1585_req
      -- CP-element group 84: 	 branch_block_stmt_1432/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1585/phi_stmt_1585_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_1432/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1585/phi_stmt_1585_sources/type_cast_1591/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_1432/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1585/phi_stmt_1585_sources/type_cast_1591/$exit
      -- 
    phi_stmt_1585_req_4636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1585_req_4636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(84), ack => phi_stmt_1585_req_1); -- 
    convTransposeA_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3912_elements(82) & convTransposeA_CP_3912_elements(83);
      gj_convTransposeA_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3912_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  output  delay-element  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	81 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (5) 
      -- CP-element group 85: 	 branch_block_stmt_1432/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1585/$exit
      -- CP-element group 85: 	 branch_block_stmt_1432/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1585/phi_stmt_1585_sources/$exit
      -- CP-element group 85: 	 branch_block_stmt_1432/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1585/phi_stmt_1585_sources/type_cast_1589_konst_delay_trans
      -- CP-element group 85: 	 branch_block_stmt_1432/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 85: 	 branch_block_stmt_1432/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1585/phi_stmt_1585_req
      -- 
    phi_stmt_1585_req_4647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1585_req_4647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(85), ack => phi_stmt_1585_req_0); -- 
    -- Element group convTransposeA_CP_3912_elements(85) is a control-delay.
    cp_element_85_delay: control_delay_element  generic map(name => " 85_delay", delay_value => 1)  port map(req => convTransposeA_CP_3912_elements(81), ack => convTransposeA_CP_3912_elements(85), clk => clk, reset =>reset);
    -- CP-element group 86:  merge  transition  place  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1432/merge_stmt_1584_PhiAck/$entry
      -- CP-element group 86: 	 branch_block_stmt_1432/merge_stmt_1584_PhiReqMerge
      -- 
    convTransposeA_CP_3912_elements(86) <= OrReduce(convTransposeA_CP_3912_elements(84) & convTransposeA_CP_3912_elements(85));
    -- CP-element group 87:  fork  transition  place  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	37 
    -- CP-element group 87: 	39 
    -- CP-element group 87: 	45 
    -- CP-element group 87: 	47 
    -- CP-element group 87: 	49 
    -- CP-element group 87: 	53 
    -- CP-element group 87: 	54 
    -- CP-element group 87: 	52 
    -- CP-element group 87: 	41 
    -- CP-element group 87: 	42 
    -- CP-element group 87: 	43 
    -- CP-element group 87: 	32 
    -- CP-element group 87: 	33 
    -- CP-element group 87: 	35 
    -- CP-element group 87:  members (51) 
      -- CP-element group 87: 	 branch_block_stmt_1432/merge_stmt_1584__exit__
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687__entry__
      -- CP-element group 87: 	 branch_block_stmt_1432/merge_stmt_1584_PhiAck/$exit
      -- CP-element group 87: 	 branch_block_stmt_1432/merge_stmt_1584_PhiAck/phi_stmt_1585_ack
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/$entry
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1613_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1613_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1613_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1613_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1613_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1613_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1627_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1627_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1627_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1634_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_final_index_sum_regn_update_start
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_final_index_sum_regn_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1633_final_index_sum_regn_Update/req
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1634_complete/$entry
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1634_complete/req
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_Update/word_access_complete/$entry
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_Update/word_access_complete/word_0/$entry
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1638_Update/word_access_complete/word_0/cr
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1643_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1643_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1643_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1643_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1643_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1643_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1657_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1657_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1657_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1664_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_final_index_sum_regn_update_start
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_final_index_sum_regn_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/array_obj_ref_1663_final_index_sum_regn_Update/req
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1664_complete/$entry
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/addr_of_1664_complete/req
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_Update/word_access_complete/$entry
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_Update/word_access_complete/word_0/$entry
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/ptr_deref_1667_Update/word_access_complete/word_0/cr
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1673_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1673_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1673_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1673_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1673_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1432/assign_stmt_1598_to_assign_stmt_1687/type_cast_1673_Update/cr
      -- 
    phi_stmt_1585_ack_4652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1585_ack_0, ack => convTransposeA_CP_3912_elements(87)); -- 
    rr_4179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(87), ack => type_cast_1613_inst_req_0); -- 
    cr_4184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(87), ack => type_cast_1613_inst_req_1); -- 
    cr_4198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(87), ack => type_cast_1627_inst_req_1); -- 
    req_4229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(87), ack => array_obj_ref_1633_index_offset_req_1); -- 
    req_4244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(87), ack => addr_of_1634_final_reg_req_1); -- 
    cr_4289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(87), ack => ptr_deref_1638_load_0_req_1); -- 
    rr_4303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(87), ack => type_cast_1643_inst_req_0); -- 
    cr_4308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(87), ack => type_cast_1643_inst_req_1); -- 
    cr_4322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(87), ack => type_cast_1657_inst_req_1); -- 
    req_4353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(87), ack => array_obj_ref_1663_index_offset_req_1); -- 
    req_4368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(87), ack => addr_of_1664_final_reg_req_1); -- 
    cr_4418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(87), ack => ptr_deref_1667_store_0_req_1); -- 
    rr_4427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(87), ack => type_cast_1673_inst_req_0); -- 
    cr_4432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3912_elements(87), ack => type_cast_1673_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1621_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1651_wire : std_logic_vector(31 downto 0);
    signal R_idxprom85_1662_resized : std_logic_vector(13 downto 0);
    signal R_idxprom85_1662_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1632_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1632_scaled : std_logic_vector(13 downto 0);
    signal add32_1603 : std_logic_vector(15 downto 0);
    signal add76_1608 : std_logic_vector(15 downto 0);
    signal add90_1680 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1633_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1633_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1633_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1633_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1633_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1633_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1663_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1663_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1663_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1663_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1663_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1663_root_address : std_logic_vector(13 downto 0);
    signal arrayidx80_1635 : std_logic_vector(31 downto 0);
    signal arrayidx86_1665 : std_logic_vector(31 downto 0);
    signal call11_1453 : std_logic_vector(15 downto 0);
    signal call13_1456 : std_logic_vector(15 downto 0);
    signal call14_1459 : std_logic_vector(15 downto 0);
    signal call15_1462 : std_logic_vector(15 downto 0);
    signal call17_1465 : std_logic_vector(15 downto 0);
    signal call19_1468 : std_logic_vector(15 downto 0);
    signal call1_1438 : std_logic_vector(15 downto 0);
    signal call3_1441 : std_logic_vector(15 downto 0);
    signal call5_1444 : std_logic_vector(15 downto 0);
    signal call7_1447 : std_logic_vector(15 downto 0);
    signal call9_1450 : std_logic_vector(15 downto 0);
    signal call_1435 : std_logic_vector(15 downto 0);
    signal cmp105_1718 : std_logic_vector(0 downto 0);
    signal cmp116_1744 : std_logic_vector(0 downto 0);
    signal cmp_1687 : std_logic_vector(0 downto 0);
    signal conv101_1713 : std_logic_vector(31 downto 0);
    signal conv104_1477 : std_logic_vector(31 downto 0);
    signal conv111_1739 : std_logic_vector(31 downto 0);
    signal conv114_1487 : std_logic_vector(31 downto 0);
    signal conv79_1614 : std_logic_vector(31 downto 0);
    signal conv83_1644 : std_logic_vector(31 downto 0);
    signal conv89_1674 : std_logic_vector(31 downto 0);
    signal conv93_1473 : std_logic_vector(31 downto 0);
    signal div115_1493 : std_logic_vector(31 downto 0);
    signal div_1483 : std_logic_vector(31 downto 0);
    signal idxprom85_1658 : std_logic_vector(63 downto 0);
    signal idxprom_1628 : std_logic_vector(63 downto 0);
    signal inc109_1722 : std_logic_vector(15 downto 0);
    signal inc109x_xinput_dim0x_x2_1727 : std_logic_vector(15 downto 0);
    signal inc_1708 : std_logic_vector(15 downto 0);
    signal indvar_1585 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_1700 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_1525 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_1518 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1734 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1598 : std_logic_vector(15 downto 0);
    signal ptr_deref_1638_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1638_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1638_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1638_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1638_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1667_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1667_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1667_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1667_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1667_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1667_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr84_1653 : std_logic_vector(31 downto 0);
    signal shr_1623 : std_logic_vector(31 downto 0);
    signal tmp10_1582 : std_logic_vector(15 downto 0);
    signal tmp143_1537 : std_logic_vector(15 downto 0);
    signal tmp144_1542 : std_logic_vector(15 downto 0);
    signal tmp145_1547 : std_logic_vector(15 downto 0);
    signal tmp1_1504 : std_logic_vector(15 downto 0);
    signal tmp2_1552 : std_logic_vector(15 downto 0);
    signal tmp3_1557 : std_logic_vector(15 downto 0);
    signal tmp4_1510 : std_logic_vector(15 downto 0);
    signal tmp5_1515 : std_logic_vector(15 downto 0);
    signal tmp6_1562 : std_logic_vector(15 downto 0);
    signal tmp7_1567 : std_logic_vector(15 downto 0);
    signal tmp81_1639 : std_logic_vector(63 downto 0);
    signal tmp8_1572 : std_logic_vector(15 downto 0);
    signal tmp9_1577 : std_logic_vector(15 downto 0);
    signal tmp_1499 : std_logic_vector(15 downto 0);
    signal type_cast_1481_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1491_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1497_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1508_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1522_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1524_wire : std_logic_vector(15 downto 0);
    signal type_cast_1529_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1531_wire : std_logic_vector(15 downto 0);
    signal type_cast_1589_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1591_wire : std_logic_vector(15 downto 0);
    signal type_cast_1596_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1612_wire : std_logic_vector(31 downto 0);
    signal type_cast_1617_wire : std_logic_vector(31 downto 0);
    signal type_cast_1620_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1626_wire : std_logic_vector(63 downto 0);
    signal type_cast_1642_wire : std_logic_vector(31 downto 0);
    signal type_cast_1647_wire : std_logic_vector(31 downto 0);
    signal type_cast_1650_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1656_wire : std_logic_vector(63 downto 0);
    signal type_cast_1672_wire : std_logic_vector(31 downto 0);
    signal type_cast_1678_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1683_wire : std_logic_vector(31 downto 0);
    signal type_cast_1685_wire : std_logic_vector(31 downto 0);
    signal type_cast_1698_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1706_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1711_wire : std_logic_vector(31 downto 0);
    signal type_cast_1731_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1737_wire : std_logic_vector(31 downto 0);
    signal type_cast_1755_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_1633_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1633_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1633_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1633_resized_base_address <= "00000000000000";
    array_obj_ref_1663_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1663_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1663_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1663_resized_base_address <= "00000000000000";
    ptr_deref_1638_word_offset_0 <= "00000000000000";
    ptr_deref_1667_word_offset_0 <= "00000000000000";
    type_cast_1481_wire_constant <= "00000000000000000000000000000001";
    type_cast_1491_wire_constant <= "00000000000000000000000000000001";
    type_cast_1497_wire_constant <= "1111111111111111";
    type_cast_1508_wire_constant <= "1111111111111111";
    type_cast_1522_wire_constant <= "0000000000000000";
    type_cast_1529_wire_constant <= "0000000000000000";
    type_cast_1589_wire_constant <= "0000000000000000";
    type_cast_1596_wire_constant <= "0000000000000100";
    type_cast_1620_wire_constant <= "00000000000000000000000000000010";
    type_cast_1650_wire_constant <= "00000000000000000000000000000010";
    type_cast_1678_wire_constant <= "00000000000000000000000000000100";
    type_cast_1698_wire_constant <= "0000000000000001";
    type_cast_1706_wire_constant <= "0000000000000001";
    type_cast_1731_wire_constant <= "0000000000000000";
    type_cast_1755_wire_constant <= "0000000000000001";
    phi_stmt_1518: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1522_wire_constant & type_cast_1524_wire;
      req <= phi_stmt_1518_req_0 & phi_stmt_1518_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1518",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1518_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_1518,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1518
    phi_stmt_1525: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1529_wire_constant & type_cast_1531_wire;
      req <= phi_stmt_1525_req_0 & phi_stmt_1525_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1525",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1525_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_1525,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1525
    phi_stmt_1585: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1589_wire_constant & type_cast_1591_wire;
      req <= phi_stmt_1585_req_0 & phi_stmt_1585_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1585",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1585_ack_0,
          idata => idata,
          odata => indvar_1585,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1585
    -- flow-through select operator MUX_1733_inst
    input_dim1x_x2_1734 <= type_cast_1731_wire_constant when (cmp105_1718(0) /=  '0') else inc_1708;
    addr_of_1634_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1634_final_reg_req_0;
      addr_of_1634_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1634_final_reg_req_1;
      addr_of_1634_final_reg_ack_1<= rack(0);
      addr_of_1634_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1634_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1633_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx80_1635,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1664_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1664_final_reg_req_0;
      addr_of_1664_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1664_final_reg_req_1;
      addr_of_1664_final_reg_ack_1<= rack(0);
      addr_of_1664_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1664_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1663_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx86_1665,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1472_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1472_inst_req_0;
      type_cast_1472_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1472_inst_req_1;
      type_cast_1472_inst_ack_1<= rack(0);
      type_cast_1472_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1472_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1441,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv93_1473,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1476_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1476_inst_req_0;
      type_cast_1476_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1476_inst_req_1;
      type_cast_1476_inst_ack_1<= rack(0);
      type_cast_1476_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1476_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_1438,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_1477,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1486_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1486_inst_req_0;
      type_cast_1486_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1486_inst_req_1;
      type_cast_1486_inst_ack_1<= rack(0);
      type_cast_1486_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1486_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1435,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv114_1487,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1524_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1524_inst_req_0;
      type_cast_1524_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1524_inst_req_1;
      type_cast_1524_inst_ack_1<= rack(0);
      type_cast_1524_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1524_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1734,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1524_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1531_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1531_inst_req_0;
      type_cast_1531_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1531_inst_req_1;
      type_cast_1531_inst_ack_1<= rack(0);
      type_cast_1531_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1531_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc109x_xinput_dim0x_x2_1727,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1531_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1591_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1591_inst_req_0;
      type_cast_1591_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1591_inst_req_1;
      type_cast_1591_inst_ack_1<= rack(0);
      type_cast_1591_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1591_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1700,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1591_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1613_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1613_inst_req_0;
      type_cast_1613_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1613_inst_req_1;
      type_cast_1613_inst_ack_1<= rack(0);
      type_cast_1613_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1613_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1612_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_1614,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1617_inst
    process(conv79_1614) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv79_1614(31 downto 0);
      type_cast_1617_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1622_inst
    process(ASHR_i32_i32_1621_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1621_wire(31 downto 0);
      shr_1623 <= tmp_var; -- 
    end process;
    type_cast_1627_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1627_inst_req_0;
      type_cast_1627_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1627_inst_req_1;
      type_cast_1627_inst_ack_1<= rack(0);
      type_cast_1627_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1627_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1626_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1628,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1643_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1643_inst_req_0;
      type_cast_1643_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1643_inst_req_1;
      type_cast_1643_inst_ack_1<= rack(0);
      type_cast_1643_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1643_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1642_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_1644,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1647_inst
    process(conv83_1644) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv83_1644(31 downto 0);
      type_cast_1647_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1652_inst
    process(ASHR_i32_i32_1651_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1651_wire(31 downto 0);
      shr84_1653 <= tmp_var; -- 
    end process;
    type_cast_1657_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1657_inst_req_0;
      type_cast_1657_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1657_inst_req_1;
      type_cast_1657_inst_ack_1<= rack(0);
      type_cast_1657_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1657_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1656_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom85_1658,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1673_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1673_inst_req_0;
      type_cast_1673_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1673_inst_req_1;
      type_cast_1673_inst_ack_1<= rack(0);
      type_cast_1673_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1673_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1672_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv89_1674,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1683_inst
    process(add90_1680) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add90_1680(31 downto 0);
      type_cast_1683_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1685_inst
    process(conv93_1473) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv93_1473(31 downto 0);
      type_cast_1685_wire <= tmp_var; -- 
    end process;
    type_cast_1712_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1712_inst_req_0;
      type_cast_1712_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1712_inst_req_1;
      type_cast_1712_inst_ack_1<= rack(0);
      type_cast_1712_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1712_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1711_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv101_1713,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1721_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1721_inst_req_0;
      type_cast_1721_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1721_inst_req_1;
      type_cast_1721_inst_ack_1<= rack(0);
      type_cast_1721_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1721_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp105_1718,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc109_1722,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1738_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1738_inst_req_0;
      type_cast_1738_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1738_inst_req_1;
      type_cast_1738_inst_ack_1<= rack(0);
      type_cast_1738_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1738_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1737_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv111_1739,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1633_index_1_rename
    process(R_idxprom_1632_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1632_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1632_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1633_index_1_resize
    process(idxprom_1628) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1628;
      ov := iv(13 downto 0);
      R_idxprom_1632_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1633_root_address_inst
    process(array_obj_ref_1633_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1633_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1633_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1663_index_1_rename
    process(R_idxprom85_1662_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom85_1662_resized;
      ov(13 downto 0) := iv;
      R_idxprom85_1662_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1663_index_1_resize
    process(idxprom85_1658) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom85_1658;
      ov := iv(13 downto 0);
      R_idxprom85_1662_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1663_root_address_inst
    process(array_obj_ref_1663_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1663_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1663_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1638_addr_0
    process(ptr_deref_1638_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1638_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1638_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1638_base_resize
    process(arrayidx80_1635) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx80_1635;
      ov := iv(13 downto 0);
      ptr_deref_1638_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1638_gather_scatter
    process(ptr_deref_1638_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1638_data_0;
      ov(63 downto 0) := iv;
      tmp81_1639 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1638_root_address_inst
    process(ptr_deref_1638_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1638_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1638_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1667_addr_0
    process(ptr_deref_1667_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1667_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1667_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1667_base_resize
    process(arrayidx86_1665) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx86_1665;
      ov := iv(13 downto 0);
      ptr_deref_1667_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1667_gather_scatter
    process(tmp81_1639) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp81_1639;
      ov(63 downto 0) := iv;
      ptr_deref_1667_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1667_root_address_inst
    process(ptr_deref_1667_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1667_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1667_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1688_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1687;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1688_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1688_branch_req_0,
          ack0 => if_stmt_1688_branch_ack_0,
          ack1 => if_stmt_1688_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1745_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp116_1744;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1745_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1745_branch_req_0,
          ack0 => if_stmt_1745_branch_ack_0,
          ack1 => if_stmt_1745_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1498_inst
    process(call9_1450) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1450, type_cast_1497_wire_constant, tmp_var);
      tmp_1499 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1509_inst
    process(call7_1447) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1447, type_cast_1508_wire_constant, tmp_var);
      tmp4_1510 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1541_inst
    process(input_dim1x_x1x_xph_1518, tmp143_1537) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1518, tmp143_1537, tmp_var);
      tmp144_1542 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1556_inst
    process(tmp1_1504, tmp2_1552) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp1_1504, tmp2_1552, tmp_var);
      tmp3_1557 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1566_inst
    process(tmp5_1515, tmp6_1562) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp5_1515, tmp6_1562, tmp_var);
      tmp7_1567 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1576_inst
    process(tmp3_1557, tmp8_1572) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_1557, tmp8_1572, tmp_var);
      tmp9_1577 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1602_inst
    process(tmp145_1547, input_dim2x_x1_1598) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp145_1547, input_dim2x_x1_1598, tmp_var);
      add32_1603 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1607_inst
    process(tmp10_1582, input_dim2x_x1_1598) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp10_1582, input_dim2x_x1_1598, tmp_var);
      add76_1608 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1699_inst
    process(indvar_1585) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1585, type_cast_1698_wire_constant, tmp_var);
      indvarx_xnext_1700 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1707_inst
    process(input_dim1x_x1x_xph_1518) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1518, type_cast_1706_wire_constant, tmp_var);
      inc_1708 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1726_inst
    process(inc109_1722, input_dim0x_x2x_xph_1525) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc109_1722, input_dim0x_x2x_xph_1525, tmp_var);
      inc109x_xinput_dim0x_x2_1727 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1679_inst
    process(conv89_1674) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv89_1674, type_cast_1678_wire_constant, tmp_var);
      add90_1680 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1621_inst
    process(type_cast_1617_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1617_wire, type_cast_1620_wire_constant, tmp_var);
      ASHR_i32_i32_1621_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1651_inst
    process(type_cast_1647_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1647_wire, type_cast_1650_wire_constant, tmp_var);
      ASHR_i32_i32_1651_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1717_inst
    process(conv101_1713, div_1483) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv101_1713, div_1483, tmp_var);
      cmp105_1718 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1743_inst
    process(conv111_1739, div115_1493) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv111_1739, div115_1493, tmp_var);
      cmp116_1744 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1482_inst
    process(conv104_1477) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv104_1477, type_cast_1481_wire_constant, tmp_var);
      div_1483 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1492_inst
    process(conv114_1487) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv114_1487, type_cast_1491_wire_constant, tmp_var);
      div115_1493 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1536_inst
    process(call1_1438, input_dim0x_x2x_xph_1525) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call1_1438, input_dim0x_x2x_xph_1525, tmp_var);
      tmp143_1537 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1546_inst
    process(call3_1441, tmp144_1542) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call3_1441, tmp144_1542, tmp_var);
      tmp145_1547 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1551_inst
    process(call13_1456, input_dim1x_x1x_xph_1518) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_1456, input_dim1x_x1x_xph_1518, tmp_var);
      tmp2_1552 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1561_inst
    process(call13_1456, input_dim0x_x2x_xph_1525) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_1456, input_dim0x_x2x_xph_1525, tmp_var);
      tmp6_1562 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1571_inst
    process(call17_1465, tmp7_1567) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call17_1465, tmp7_1567, tmp_var);
      tmp8_1572 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1581_inst
    process(call19_1468, tmp9_1577) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call19_1468, tmp9_1577, tmp_var);
      tmp10_1582 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1597_inst
    process(indvar_1585) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1585, type_cast_1596_wire_constant, tmp_var);
      input_dim2x_x1_1598 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1686_inst
    process(type_cast_1683_wire, type_cast_1685_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1683_wire, type_cast_1685_wire, tmp_var);
      cmp_1687 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1503_inst
    process(tmp_1499, call14_1459) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp_1499, call14_1459, tmp_var);
      tmp1_1504 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1514_inst
    process(tmp4_1510, call14_1459) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp4_1510, call14_1459, tmp_var);
      tmp5_1515 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_1633_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1632_scaled;
      array_obj_ref_1633_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1633_index_offset_req_0;
      array_obj_ref_1633_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1633_index_offset_req_1;
      array_obj_ref_1633_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_1663_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom85_1662_scaled;
      array_obj_ref_1663_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1663_index_offset_req_0;
      array_obj_ref_1663_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1663_index_offset_req_1;
      array_obj_ref_1663_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- unary operator type_cast_1612_inst
    process(add32_1603) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add32_1603, tmp_var);
      type_cast_1612_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1626_inst
    process(shr_1623) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1623, tmp_var);
      type_cast_1626_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1642_inst
    process(add76_1608) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add76_1608, tmp_var);
      type_cast_1642_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1656_inst
    process(shr84_1653) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr84_1653, tmp_var);
      type_cast_1656_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1672_inst
    process(input_dim2x_x1_1598) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_1598, tmp_var);
      type_cast_1672_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1711_inst
    process(inc_1708) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_1708, tmp_var);
      type_cast_1711_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1737_inst
    process(inc109x_xinput_dim0x_x2_1727) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc109x_xinput_dim0x_x2_1727, tmp_var);
      type_cast_1737_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1638_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1638_load_0_req_0;
      ptr_deref_1638_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1638_load_0_req_1;
      ptr_deref_1638_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1638_word_address_0;
      ptr_deref_1638_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1667_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1667_store_0_req_0;
      ptr_deref_1667_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1667_store_0_req_1;
      ptr_deref_1667_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1667_word_address_0;
      data_in <= ptr_deref_1667_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1437_inst RPIPE_Block0_start_1452_inst RPIPE_Block0_start_1458_inst RPIPE_Block0_start_1455_inst RPIPE_Block0_start_1449_inst RPIPE_Block0_start_1440_inst RPIPE_Block0_start_1443_inst RPIPE_Block0_start_1446_inst RPIPE_Block0_start_1461_inst RPIPE_Block0_start_1434_inst RPIPE_Block0_start_1464_inst RPIPE_Block0_start_1467_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(191 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 11 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 11 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant outBUFs : IntegerArray(11 downto 0) := (11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      reqL_unguarded(11) <= RPIPE_Block0_start_1437_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block0_start_1452_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block0_start_1458_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block0_start_1455_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block0_start_1449_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block0_start_1440_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block0_start_1443_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block0_start_1446_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block0_start_1461_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block0_start_1434_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block0_start_1464_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block0_start_1467_inst_req_0;
      RPIPE_Block0_start_1437_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block0_start_1452_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block0_start_1458_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block0_start_1455_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block0_start_1449_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block0_start_1440_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block0_start_1443_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block0_start_1446_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block0_start_1461_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block0_start_1434_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block0_start_1464_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block0_start_1467_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(11) <= RPIPE_Block0_start_1437_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block0_start_1452_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block0_start_1458_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block0_start_1455_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block0_start_1449_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block0_start_1440_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block0_start_1443_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block0_start_1446_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block0_start_1461_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block0_start_1434_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block0_start_1464_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block0_start_1467_inst_req_1;
      RPIPE_Block0_start_1437_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block0_start_1452_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block0_start_1458_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block0_start_1455_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block0_start_1449_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block0_start_1440_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block0_start_1443_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block0_start_1446_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block0_start_1461_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block0_start_1434_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block0_start_1464_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block0_start_1467_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      call1_1438 <= data_out(191 downto 176);
      call11_1453 <= data_out(175 downto 160);
      call14_1459 <= data_out(159 downto 144);
      call13_1456 <= data_out(143 downto 128);
      call9_1450 <= data_out(127 downto 112);
      call3_1441 <= data_out(111 downto 96);
      call5_1444 <= data_out(95 downto 80);
      call7_1447 <= data_out(79 downto 64);
      call15_1462 <= data_out(63 downto 48);
      call_1435 <= data_out(47 downto 32);
      call17_1465 <= data_out(31 downto 16);
      call19_1468 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 12,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1753_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1753_inst_req_0;
      WPIPE_Block0_done_1753_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1753_inst_req_1;
      WPIPE_Block0_done_1753_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1755_wire_constant;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_4693_start: Boolean;
  signal convTransposeB_CP_4693_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block1_start_1797_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1773_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1785_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1776_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1785_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1794_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1776_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1770_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1764_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1794_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1794_inst_req_0 : boolean;
  signal type_cast_1812_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1797_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1782_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1785_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1770_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1785_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1791_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1770_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1773_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1782_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1767_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1782_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1767_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1791_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1764_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1764_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1791_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1767_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1779_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1767_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1779_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1779_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1791_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1776_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1776_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1782_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1779_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1770_inst_req_0 : boolean;
  signal type_cast_1812_inst_ack_0 : boolean;
  signal type_cast_1808_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1764_inst_req_1 : boolean;
  signal type_cast_1816_inst_req_0 : boolean;
  signal type_cast_1816_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1788_inst_ack_1 : boolean;
  signal type_cast_1812_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1788_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1797_inst_ack_1 : boolean;
  signal type_cast_1812_inst_ack_1 : boolean;
  signal array_obj_ref_1961_index_offset_req_1 : boolean;
  signal array_obj_ref_1961_index_offset_ack_1 : boolean;
  signal type_cast_1808_inst_req_1 : boolean;
  signal type_cast_1808_inst_ack_0 : boolean;
  signal type_cast_1808_inst_req_0 : boolean;
  signal type_cast_1955_inst_req_1 : boolean;
  signal type_cast_1955_inst_ack_1 : boolean;
  signal array_obj_ref_1961_index_offset_ack_0 : boolean;
  signal array_obj_ref_1961_index_offset_req_0 : boolean;
  signal type_cast_1941_inst_req_1 : boolean;
  signal type_cast_1941_inst_ack_1 : boolean;
  signal type_cast_1941_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1773_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1788_inst_ack_0 : boolean;
  signal addr_of_1962_final_reg_req_1 : boolean;
  signal addr_of_1962_final_reg_ack_1 : boolean;
  signal RPIPE_Block1_start_1773_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1797_inst_req_1 : boolean;
  signal addr_of_1962_final_reg_req_0 : boolean;
  signal addr_of_1962_final_reg_ack_0 : boolean;
  signal type_cast_1816_inst_req_1 : boolean;
  signal type_cast_1816_inst_ack_1 : boolean;
  signal type_cast_1941_inst_req_0 : boolean;
  signal type_cast_1955_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1788_inst_req_0 : boolean;
  signal type_cast_1955_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1794_inst_ack_0 : boolean;
  signal ptr_deref_1966_load_0_req_0 : boolean;
  signal ptr_deref_1966_load_0_ack_0 : boolean;
  signal ptr_deref_1966_load_0_req_1 : boolean;
  signal ptr_deref_1966_load_0_ack_1 : boolean;
  signal type_cast_1971_inst_req_0 : boolean;
  signal type_cast_1971_inst_ack_0 : boolean;
  signal type_cast_1971_inst_req_1 : boolean;
  signal type_cast_1971_inst_ack_1 : boolean;
  signal type_cast_1985_inst_req_0 : boolean;
  signal type_cast_1985_inst_ack_0 : boolean;
  signal type_cast_1985_inst_req_1 : boolean;
  signal type_cast_1985_inst_ack_1 : boolean;
  signal array_obj_ref_1991_index_offset_req_0 : boolean;
  signal array_obj_ref_1991_index_offset_ack_0 : boolean;
  signal array_obj_ref_1991_index_offset_req_1 : boolean;
  signal array_obj_ref_1991_index_offset_ack_1 : boolean;
  signal addr_of_1992_final_reg_req_0 : boolean;
  signal addr_of_1992_final_reg_ack_0 : boolean;
  signal addr_of_1992_final_reg_req_1 : boolean;
  signal addr_of_1992_final_reg_ack_1 : boolean;
  signal ptr_deref_1995_store_0_req_0 : boolean;
  signal ptr_deref_1995_store_0_ack_0 : boolean;
  signal ptr_deref_1995_store_0_req_1 : boolean;
  signal ptr_deref_1995_store_0_ack_1 : boolean;
  signal type_cast_2001_inst_req_0 : boolean;
  signal type_cast_2001_inst_ack_0 : boolean;
  signal type_cast_2001_inst_req_1 : boolean;
  signal type_cast_2001_inst_ack_1 : boolean;
  signal if_stmt_2016_branch_req_0 : boolean;
  signal if_stmt_2016_branch_ack_1 : boolean;
  signal if_stmt_2016_branch_ack_0 : boolean;
  signal type_cast_2040_inst_req_0 : boolean;
  signal type_cast_2040_inst_ack_0 : boolean;
  signal type_cast_2040_inst_req_1 : boolean;
  signal type_cast_2040_inst_ack_1 : boolean;
  signal type_cast_2055_inst_req_0 : boolean;
  signal type_cast_2055_inst_ack_0 : boolean;
  signal type_cast_2055_inst_req_1 : boolean;
  signal type_cast_2055_inst_ack_1 : boolean;
  signal type_cast_2065_inst_req_0 : boolean;
  signal type_cast_2065_inst_ack_0 : boolean;
  signal type_cast_2065_inst_req_1 : boolean;
  signal type_cast_2065_inst_ack_1 : boolean;
  signal if_stmt_2072_branch_req_0 : boolean;
  signal if_stmt_2072_branch_ack_1 : boolean;
  signal if_stmt_2072_branch_ack_0 : boolean;
  signal WPIPE_Block1_done_2080_inst_req_0 : boolean;
  signal WPIPE_Block1_done_2080_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_2080_inst_req_1 : boolean;
  signal WPIPE_Block1_done_2080_inst_ack_1 : boolean;
  signal type_cast_1851_inst_req_0 : boolean;
  signal type_cast_1851_inst_ack_0 : boolean;
  signal type_cast_1851_inst_req_1 : boolean;
  signal type_cast_1851_inst_ack_1 : boolean;
  signal phi_stmt_1848_req_0 : boolean;
  signal phi_stmt_1854_req_0 : boolean;
  signal type_cast_1853_inst_req_0 : boolean;
  signal type_cast_1853_inst_ack_0 : boolean;
  signal type_cast_1853_inst_req_1 : boolean;
  signal type_cast_1853_inst_ack_1 : boolean;
  signal phi_stmt_1848_req_1 : boolean;
  signal type_cast_1860_inst_req_0 : boolean;
  signal type_cast_1860_inst_ack_0 : boolean;
  signal type_cast_1860_inst_req_1 : boolean;
  signal type_cast_1860_inst_ack_1 : boolean;
  signal phi_stmt_1854_req_1 : boolean;
  signal phi_stmt_1848_ack_0 : boolean;
  signal phi_stmt_1854_ack_0 : boolean;
  signal type_cast_1917_inst_req_0 : boolean;
  signal type_cast_1917_inst_ack_0 : boolean;
  signal type_cast_1917_inst_req_1 : boolean;
  signal type_cast_1917_inst_ack_1 : boolean;
  signal phi_stmt_1914_req_0 : boolean;
  signal phi_stmt_1914_req_1 : boolean;
  signal phi_stmt_1914_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_4693_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4693_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_4693_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4693_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_4693: Block -- control-path 
    signal convTransposeB_CP_4693_elements: BooleanArray(89 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_4693_elements(0) <= convTransposeB_CP_4693_start;
    convTransposeB_CP_4693_symbol <= convTransposeB_CP_4693_elements(67);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798__entry__
      -- CP-element group 0: 	 branch_block_stmt_1762/branch_block_stmt_1762__entry__
      -- CP-element group 0: 	 branch_block_stmt_1762/$entry
      -- CP-element group 0: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1764_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1764_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/$entry
      -- CP-element group 0: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1764_sample_start_
      -- 
    rr_4741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(0), ack => RPIPE_Block1_start_1764_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1764_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1764_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1764_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1764_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1764_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1764_update_start_
      -- 
    ra_4742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1764_inst_ack_0, ack => convTransposeB_CP_4693_elements(1)); -- 
    cr_4746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(1), ack => RPIPE_Block1_start_1764_inst_req_1); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1767_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1764_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1764_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1767_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1767_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1764_Update/$exit
      -- 
    ca_4747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1764_inst_ack_1, ack => convTransposeB_CP_4693_elements(2)); -- 
    rr_4755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(2), ack => RPIPE_Block1_start_1767_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1767_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1767_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1767_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1767_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1767_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1767_Update/cr
      -- 
    ra_4756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1767_inst_ack_0, ack => convTransposeB_CP_4693_elements(3)); -- 
    cr_4760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(3), ack => RPIPE_Block1_start_1767_inst_req_1); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1767_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1767_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1767_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1770_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1770_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1770_Sample/rr
      -- 
    ca_4761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1767_inst_ack_1, ack => convTransposeB_CP_4693_elements(4)); -- 
    rr_4769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(4), ack => RPIPE_Block1_start_1770_inst_req_0); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1770_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1770_Update/cr
      -- CP-element group 5: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1770_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1770_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1770_update_start_
      -- CP-element group 5: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1770_Sample/$exit
      -- 
    ra_4770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1770_inst_ack_0, ack => convTransposeB_CP_4693_elements(5)); -- 
    cr_4774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(5), ack => RPIPE_Block1_start_1770_inst_req_1); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1770_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1770_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1773_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1770_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1773_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1773_Sample/$entry
      -- 
    ca_4775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1770_inst_ack_1, ack => convTransposeB_CP_4693_elements(6)); -- 
    rr_4783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(6), ack => RPIPE_Block1_start_1773_inst_req_0); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1773_Update/cr
      -- CP-element group 7: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1773_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1773_update_start_
      -- CP-element group 7: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1773_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1773_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1773_Sample/$exit
      -- 
    ra_4784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1773_inst_ack_0, ack => convTransposeB_CP_4693_elements(7)); -- 
    cr_4788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(7), ack => RPIPE_Block1_start_1773_inst_req_1); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1773_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1776_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1776_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1776_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1773_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1773_update_completed_
      -- 
    ca_4789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1773_inst_ack_1, ack => convTransposeB_CP_4693_elements(8)); -- 
    rr_4797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(8), ack => RPIPE_Block1_start_1776_inst_req_0); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1776_Update/cr
      -- CP-element group 9: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1776_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1776_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1776_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1776_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1776_Update/$entry
      -- 
    ra_4798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1776_inst_ack_0, ack => convTransposeB_CP_4693_elements(9)); -- 
    cr_4802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(9), ack => RPIPE_Block1_start_1776_inst_req_1); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1776_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1779_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1779_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1776_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1779_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1776_Update/$exit
      -- 
    ca_4803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1776_inst_ack_1, ack => convTransposeB_CP_4693_elements(10)); -- 
    rr_4811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(10), ack => RPIPE_Block1_start_1779_inst_req_0); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1779_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1779_update_start_
      -- CP-element group 11: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1779_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1779_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1779_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1779_Update/cr
      -- 
    ra_4812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1779_inst_ack_0, ack => convTransposeB_CP_4693_elements(11)); -- 
    cr_4816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(11), ack => RPIPE_Block1_start_1779_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1779_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1782_Sample/rr
      -- CP-element group 12: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1779_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1779_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1782_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1782_sample_start_
      -- 
    ca_4817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1779_inst_ack_1, ack => convTransposeB_CP_4693_elements(12)); -- 
    rr_4825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(12), ack => RPIPE_Block1_start_1782_inst_req_0); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1782_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1782_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1782_Update/cr
      -- CP-element group 13: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1782_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1782_update_start_
      -- CP-element group 13: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1782_sample_completed_
      -- 
    ra_4826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1782_inst_ack_0, ack => convTransposeB_CP_4693_elements(13)); -- 
    cr_4830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(13), ack => RPIPE_Block1_start_1782_inst_req_1); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1785_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1785_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1782_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1782_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1782_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1785_sample_start_
      -- 
    ca_4831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1782_inst_ack_1, ack => convTransposeB_CP_4693_elements(14)); -- 
    rr_4839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(14), ack => RPIPE_Block1_start_1785_inst_req_0); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1785_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1785_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1785_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1785_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1785_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1785_sample_completed_
      -- 
    ra_4840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1785_inst_ack_0, ack => convTransposeB_CP_4693_elements(15)); -- 
    cr_4844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(15), ack => RPIPE_Block1_start_1785_inst_req_1); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1785_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1785_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1788_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1785_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1788_Sample/rr
      -- CP-element group 16: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1788_Sample/$entry
      -- 
    ca_4845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1785_inst_ack_1, ack => convTransposeB_CP_4693_elements(16)); -- 
    rr_4853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(16), ack => RPIPE_Block1_start_1788_inst_req_0); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1788_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1788_update_start_
      -- CP-element group 17: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1788_Update/cr
      -- CP-element group 17: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1788_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1788_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1788_Sample/$exit
      -- 
    ra_4854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1788_inst_ack_0, ack => convTransposeB_CP_4693_elements(17)); -- 
    cr_4858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(17), ack => RPIPE_Block1_start_1788_inst_req_1); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1791_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1791_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1788_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1791_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1788_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1788_Update/$exit
      -- 
    ca_4859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1788_inst_ack_1, ack => convTransposeB_CP_4693_elements(18)); -- 
    rr_4867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(18), ack => RPIPE_Block1_start_1791_inst_req_0); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1791_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1791_update_start_
      -- CP-element group 19: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1791_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1791_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1791_Update/cr
      -- CP-element group 19: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1791_Sample/ra
      -- 
    ra_4868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1791_inst_ack_0, ack => convTransposeB_CP_4693_elements(19)); -- 
    cr_4872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(19), ack => RPIPE_Block1_start_1791_inst_req_1); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1791_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1794_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1791_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1791_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1794_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1794_Sample/$entry
      -- 
    ca_4873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1791_inst_ack_1, ack => convTransposeB_CP_4693_elements(20)); -- 
    rr_4881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(20), ack => RPIPE_Block1_start_1794_inst_req_0); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1794_Update/cr
      -- CP-element group 21: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1794_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1794_update_start_
      -- CP-element group 21: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1794_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1794_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1794_Update/$entry
      -- 
    ra_4882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1794_inst_ack_0, ack => convTransposeB_CP_4693_elements(21)); -- 
    cr_4886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(21), ack => RPIPE_Block1_start_1794_inst_req_1); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1797_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1797_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1794_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1797_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1794_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1794_update_completed_
      -- 
    ca_4887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1794_inst_ack_1, ack => convTransposeB_CP_4693_elements(22)); -- 
    rr_4895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(22), ack => RPIPE_Block1_start_1797_inst_req_0); -- 
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1797_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1797_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1797_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1797_update_start_
      -- CP-element group 23: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1797_Update/cr
      -- CP-element group 23: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1797_Update/$entry
      -- 
    ra_4896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1797_inst_ack_0, ack => convTransposeB_CP_4693_elements(23)); -- 
    cr_4900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(23), ack => RPIPE_Block1_start_1797_inst_req_1); -- 
    -- CP-element group 24:  fork  transition  place  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	30 
    -- CP-element group 24: 	25 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	27 
    -- CP-element group 24: 	28 
    -- CP-element group 24: 	29 
    -- CP-element group 24:  members (25) 
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845__entry__
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798__exit__
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1816_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1812_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1812_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/$exit
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1816_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1812_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/$entry
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1816_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1812_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1812_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1797_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1808_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1808_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1808_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1808_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1808_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1808_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1816_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1816_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1797_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1765_to_assign_stmt_1798/RPIPE_Block1_start_1797_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1816_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1812_Sample/$entry
      -- 
    ca_4901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1797_inst_ack_1, ack => convTransposeB_CP_4693_elements(24)); -- 
    rr_4926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(24), ack => type_cast_1812_inst_req_0); -- 
    rr_4940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(24), ack => type_cast_1816_inst_req_0); -- 
    cr_4931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(24), ack => type_cast_1812_inst_req_1); -- 
    cr_4917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(24), ack => type_cast_1808_inst_req_1); -- 
    rr_4912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(24), ack => type_cast_1808_inst_req_0); -- 
    cr_4945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(24), ack => type_cast_1816_inst_req_1); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1808_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1808_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1808_sample_completed_
      -- 
    ra_4913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1808_inst_ack_0, ack => convTransposeB_CP_4693_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1808_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1808_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1808_update_completed_
      -- 
    ca_4918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1808_inst_ack_1, ack => convTransposeB_CP_4693_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	24 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1812_Sample/ra
      -- CP-element group 27: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1812_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1812_sample_completed_
      -- 
    ra_4927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1812_inst_ack_0, ack => convTransposeB_CP_4693_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	24 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1812_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1812_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1812_Update/ca
      -- 
    ca_4932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1812_inst_ack_1, ack => convTransposeB_CP_4693_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	24 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1816_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1816_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1816_sample_completed_
      -- 
    ra_4941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1816_inst_ack_0, ack => convTransposeB_CP_4693_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	24 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1816_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1816_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/type_cast_1816_Update/ca
      -- 
    ca_4946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1816_inst_ack_1, ack => convTransposeB_CP_4693_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	28 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	68 
    -- CP-element group 31: 	69 
    -- CP-element group 31: 	71 
    -- CP-element group 31:  members (14) 
      -- CP-element group 31: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845__exit__
      -- CP-element group 31: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_1762/assign_stmt_1805_to_assign_stmt_1845/$exit
      -- CP-element group 31: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/$entry
      -- CP-element group 31: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1851/$entry
      -- CP-element group 31: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1851/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1851/SplitProtocol/Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1851/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1851/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1851/SplitProtocol/Update/cr
      -- CP-element group 31: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/$entry
      -- CP-element group 31: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/$entry
      -- 
    rr_5336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(31), ack => type_cast_1851_inst_req_0); -- 
    cr_5341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(31), ack => type_cast_1851_inst_req_1); -- 
    convTransposeB_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4693_elements(30) & convTransposeB_CP_4693_elements(26) & convTransposeB_CP_4693_elements(28);
      gj_convTransposeB_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4693_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	89 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1941_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1941_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1941_sample_completed_
      -- 
    ra_4961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1941_inst_ack_0, ack => convTransposeB_CP_4693_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	89 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1955_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1941_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1941_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1941_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1955_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1955_Sample/rr
      -- 
    ca_4966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1941_inst_ack_1, ack => convTransposeB_CP_4693_elements(33)); -- 
    rr_4974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(33), ack => type_cast_1955_inst_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1955_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1955_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1955_Sample/$exit
      -- 
    ra_4975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1955_inst_ack_0, ack => convTransposeB_CP_4693_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	89 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (16) 
      -- CP-element group 35: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_index_scale_1/scale_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_index_scale_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_index_scale_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_index_scale_1/scale_rename_req
      -- CP-element group 35: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_index_resize_1/index_resize_ack
      -- CP-element group 35: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_index_resize_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_index_resize_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_index_resize_1/index_resize_req
      -- CP-element group 35: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_index_resized_1
      -- CP-element group 35: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_index_scaled_1
      -- CP-element group 35: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_index_computed_1
      -- CP-element group 35: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1955_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_final_index_sum_regn_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_final_index_sum_regn_Sample/req
      -- CP-element group 35: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1955_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1955_update_completed_
      -- 
    ca_4980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1955_inst_ack_1, ack => convTransposeB_CP_4693_elements(35)); -- 
    req_5005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(35), ack => array_obj_ref_1961_index_offset_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	55 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_final_index_sum_regn_sample_complete
      -- CP-element group 36: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_final_index_sum_regn_Sample/ack
      -- CP-element group 36: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_final_index_sum_regn_Sample/$exit
      -- 
    ack_5006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1961_index_offset_ack_0, ack => convTransposeB_CP_4693_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	89 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (11) 
      -- CP-element group 37: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_final_index_sum_regn_Update/ack
      -- CP-element group 37: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_offset_calculated
      -- CP-element group 37: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1962_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_final_index_sum_regn_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1962_request/$entry
      -- CP-element group 37: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1962_request/req
      -- CP-element group 37: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_base_plus_offset/$entry
      -- CP-element group 37: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_base_plus_offset/$exit
      -- CP-element group 37: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_base_plus_offset/sum_rename_req
      -- 
    ack_5011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1961_index_offset_ack_1, ack => convTransposeB_CP_4693_elements(37)); -- 
    req_5020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(37), ack => addr_of_1962_final_reg_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1962_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1962_request/$exit
      -- CP-element group 38: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1962_request/ack
      -- 
    ack_5021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1962_final_reg_ack_0, ack => convTransposeB_CP_4693_elements(38)); -- 
    -- CP-element group 39:  join  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	89 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (24) 
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1962_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1962_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1962_complete/ack
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_base_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_word_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_base_address_resized
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_base_addr_resize/$entry
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_base_addr_resize/$exit
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_base_addr_resize/base_resize_req
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_base_addr_resize/base_resize_ack
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_word_addrgen/$entry
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_word_addrgen/$exit
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_word_addrgen/root_register_req
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_word_addrgen/root_register_ack
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_Sample/word_access_start/$entry
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_Sample/word_access_start/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_Sample/word_access_start/word_0/rr
      -- 
    ack_5026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1962_final_reg_ack_1, ack => convTransposeB_CP_4693_elements(39)); -- 
    rr_5059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(39), ack => ptr_deref_1966_load_0_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_Sample/word_access_start/$exit
      -- CP-element group 40: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_Sample/word_access_start/word_0/$exit
      -- CP-element group 40: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_Sample/word_access_start/word_0/ra
      -- 
    ra_5060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1966_load_0_ack_0, ack => convTransposeB_CP_4693_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	89 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	50 
    -- CP-element group 41:  members (9) 
      -- CP-element group 41: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_Update/word_access_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_Update/word_access_complete/word_0/$exit
      -- CP-element group 41: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_Update/word_access_complete/word_0/ca
      -- CP-element group 41: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_Update/ptr_deref_1966_Merge/$entry
      -- CP-element group 41: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_Update/ptr_deref_1966_Merge/$exit
      -- CP-element group 41: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_Update/ptr_deref_1966_Merge/merge_req
      -- CP-element group 41: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_Update/ptr_deref_1966_Merge/merge_ack
      -- 
    ca_5071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1966_load_0_ack_1, ack => convTransposeB_CP_4693_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	89 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1971_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1971_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1971_Sample/ra
      -- 
    ra_5085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1971_inst_ack_0, ack => convTransposeB_CP_4693_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	89 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1971_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1971_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1971_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1985_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1985_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1985_Sample/rr
      -- 
    ca_5090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1971_inst_ack_1, ack => convTransposeB_CP_4693_elements(43)); -- 
    rr_5098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(43), ack => type_cast_1985_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1985_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1985_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1985_Sample/ra
      -- 
    ra_5099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1985_inst_ack_0, ack => convTransposeB_CP_4693_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	89 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (16) 
      -- CP-element group 45: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_index_scale_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1985_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1985_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1985_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_index_resized_1
      -- CP-element group 45: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_index_scaled_1
      -- CP-element group 45: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_index_computed_1
      -- CP-element group 45: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_index_resize_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_index_resize_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_index_resize_1/index_resize_req
      -- CP-element group 45: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_index_resize_1/index_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_index_scale_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_index_scale_1/scale_rename_req
      -- CP-element group 45: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_index_scale_1/scale_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_final_index_sum_regn_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_final_index_sum_regn_Sample/req
      -- 
    ca_5104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1985_inst_ack_1, ack => convTransposeB_CP_4693_elements(45)); -- 
    req_5129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(45), ack => array_obj_ref_1991_index_offset_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	55 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_final_index_sum_regn_sample_complete
      -- CP-element group 46: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_final_index_sum_regn_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_final_index_sum_regn_Sample/ack
      -- 
    ack_5130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1991_index_offset_ack_0, ack => convTransposeB_CP_4693_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	89 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (11) 
      -- CP-element group 47: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1992_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_root_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_offset_calculated
      -- CP-element group 47: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_final_index_sum_regn_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_final_index_sum_regn_Update/ack
      -- CP-element group 47: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_base_plus_offset/$entry
      -- CP-element group 47: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_base_plus_offset/$exit
      -- CP-element group 47: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_base_plus_offset/sum_rename_req
      -- CP-element group 47: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_base_plus_offset/sum_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1992_request/$entry
      -- CP-element group 47: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1992_request/req
      -- 
    ack_5135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1991_index_offset_ack_1, ack => convTransposeB_CP_4693_elements(47)); -- 
    req_5144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(47), ack => addr_of_1992_final_reg_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1992_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1992_request/$exit
      -- CP-element group 48: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1992_request/ack
      -- 
    ack_5145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1992_final_reg_ack_0, ack => convTransposeB_CP_4693_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	89 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (19) 
      -- CP-element group 49: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1992_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1992_complete/$exit
      -- CP-element group 49: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1992_complete/ack
      -- CP-element group 49: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_base_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_word_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_base_address_resized
      -- CP-element group 49: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_base_addr_resize/$entry
      -- CP-element group 49: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_base_addr_resize/$exit
      -- CP-element group 49: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_base_addr_resize/base_resize_req
      -- CP-element group 49: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_base_addr_resize/base_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_word_addrgen/$entry
      -- CP-element group 49: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_word_addrgen/$exit
      -- CP-element group 49: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_word_addrgen/root_register_req
      -- CP-element group 49: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_word_addrgen/root_register_ack
      -- 
    ack_5150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1992_final_reg_ack_1, ack => convTransposeB_CP_4693_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	41 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_Sample/ptr_deref_1995_Split/$entry
      -- CP-element group 50: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_Sample/ptr_deref_1995_Split/$exit
      -- CP-element group 50: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_Sample/ptr_deref_1995_Split/split_req
      -- CP-element group 50: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_Sample/ptr_deref_1995_Split/split_ack
      -- CP-element group 50: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_Sample/word_access_start/$entry
      -- CP-element group 50: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_Sample/word_access_start/word_0/$entry
      -- CP-element group 50: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_Sample/word_access_start/word_0/rr
      -- 
    rr_5188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(50), ack => ptr_deref_1995_store_0_req_0); -- 
    convTransposeB_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4693_elements(41) & convTransposeB_CP_4693_elements(49);
      gj_convTransposeB_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4693_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_Sample/word_access_start/$exit
      -- CP-element group 51: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_Sample/word_access_start/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_Sample/word_access_start/word_0/ra
      -- 
    ra_5189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1995_store_0_ack_0, ack => convTransposeB_CP_4693_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	89 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_Update/word_access_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_Update/word_access_complete/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_Update/word_access_complete/word_0/ca
      -- 
    ca_5200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1995_store_0_ack_1, ack => convTransposeB_CP_4693_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	89 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_2001_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_2001_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_2001_Sample/ra
      -- 
    ra_5209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2001_inst_ack_0, ack => convTransposeB_CP_4693_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	89 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_2001_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_2001_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_2001_Update/ca
      -- 
    ca_5214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2001_inst_ack_1, ack => convTransposeB_CP_4693_elements(54)); -- 
    -- CP-element group 55:  branch  join  transition  place  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	36 
    -- CP-element group 55: 	52 
    -- CP-element group 55: 	54 
    -- CP-element group 55: 	46 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (10) 
      -- CP-element group 55: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015__exit__
      -- CP-element group 55: 	 branch_block_stmt_1762/if_stmt_2016__entry__
      -- CP-element group 55: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/$exit
      -- CP-element group 55: 	 branch_block_stmt_1762/if_stmt_2016_dead_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_1762/if_stmt_2016_eval_test/$entry
      -- CP-element group 55: 	 branch_block_stmt_1762/if_stmt_2016_eval_test/$exit
      -- CP-element group 55: 	 branch_block_stmt_1762/if_stmt_2016_eval_test/branch_req
      -- CP-element group 55: 	 branch_block_stmt_1762/R_cmp_2017_place
      -- CP-element group 55: 	 branch_block_stmt_1762/if_stmt_2016_if_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_1762/if_stmt_2016_else_link/$entry
      -- 
    branch_req_5222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(55), ack => if_stmt_2016_branch_req_0); -- 
    convTransposeB_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4693_elements(36) & convTransposeB_CP_4693_elements(52) & convTransposeB_CP_4693_elements(54) & convTransposeB_CP_4693_elements(46);
      gj_convTransposeB_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4693_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	84 
    -- CP-element group 56: 	85 
    -- CP-element group 56:  members (24) 
      -- CP-element group 56: 	 branch_block_stmt_1762/assign_stmt_2028__entry__
      -- CP-element group 56: 	 branch_block_stmt_1762/ifx_xthen_whilex_xbody
      -- CP-element group 56: 	 branch_block_stmt_1762/assign_stmt_2028__exit__
      -- CP-element group 56: 	 branch_block_stmt_1762/merge_stmt_2022__exit__
      -- CP-element group 56: 	 branch_block_stmt_1762/if_stmt_2016_if_link/$exit
      -- CP-element group 56: 	 branch_block_stmt_1762/if_stmt_2016_if_link/if_choice_transition
      -- CP-element group 56: 	 branch_block_stmt_1762/whilex_xbody_ifx_xthen
      -- CP-element group 56: 	 branch_block_stmt_1762/assign_stmt_2028/$entry
      -- CP-element group 56: 	 branch_block_stmt_1762/assign_stmt_2028/$exit
      -- CP-element group 56: 	 branch_block_stmt_1762/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_1762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1914/$entry
      -- CP-element group 56: 	 branch_block_stmt_1762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/$entry
      -- CP-element group 56: 	 branch_block_stmt_1762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/type_cast_1917/$entry
      -- CP-element group 56: 	 branch_block_stmt_1762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/type_cast_1917/SplitProtocol/$entry
      -- CP-element group 56: 	 branch_block_stmt_1762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/type_cast_1917/SplitProtocol/Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_1762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/type_cast_1917/SplitProtocol/Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_1762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/type_cast_1917/SplitProtocol/Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_1762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/type_cast_1917/SplitProtocol/Update/cr
      -- CP-element group 56: 	 branch_block_stmt_1762/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_1762/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_1762/merge_stmt_2022_PhiReqMerge
      -- CP-element group 56: 	 branch_block_stmt_1762/merge_stmt_2022_PhiAck/$entry
      -- CP-element group 56: 	 branch_block_stmt_1762/merge_stmt_2022_PhiAck/$exit
      -- CP-element group 56: 	 branch_block_stmt_1762/merge_stmt_2022_PhiAck/dummy
      -- 
    if_choice_transition_5227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2016_branch_ack_1, ack => convTransposeB_CP_4693_elements(56)); -- 
    rr_5425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(56), ack => type_cast_1917_inst_req_0); -- 
    cr_5430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(56), ack => type_cast_1917_inst_req_1); -- 
    -- CP-element group 57:  fork  transition  place  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	59 
    -- CP-element group 57: 	61 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (24) 
      -- CP-element group 57: 	 branch_block_stmt_1762/merge_stmt_2030__exit__
      -- CP-element group 57: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071__entry__
      -- CP-element group 57: 	 branch_block_stmt_1762/if_stmt_2016_else_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_1762/if_stmt_2016_else_link/else_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_1762/whilex_xbody_ifx_xelse
      -- CP-element group 57: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/$entry
      -- CP-element group 57: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2040_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2040_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2040_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2040_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2040_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2040_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2055_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2055_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2055_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2065_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2065_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2065_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1762/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_1762/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_1762/merge_stmt_2030_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_1762/merge_stmt_2030_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_1762/merge_stmt_2030_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_1762/merge_stmt_2030_PhiAck/dummy
      -- 
    else_choice_transition_5231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2016_branch_ack_0, ack => convTransposeB_CP_4693_elements(57)); -- 
    rr_5247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(57), ack => type_cast_2040_inst_req_0); -- 
    cr_5252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(57), ack => type_cast_2040_inst_req_1); -- 
    cr_5266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(57), ack => type_cast_2055_inst_req_1); -- 
    cr_5280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(57), ack => type_cast_2065_inst_req_1); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2040_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2040_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2040_Sample/ra
      -- 
    ra_5248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2040_inst_ack_0, ack => convTransposeB_CP_4693_elements(58)); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2040_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2040_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2040_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2055_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2055_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2055_Sample/rr
      -- 
    ca_5253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2040_inst_ack_1, ack => convTransposeB_CP_4693_elements(59)); -- 
    rr_5261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(59), ack => type_cast_2055_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2055_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2055_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2055_Sample/ra
      -- 
    ra_5262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2055_inst_ack_0, ack => convTransposeB_CP_4693_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	57 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2055_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2055_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2055_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2065_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2065_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2065_Sample/rr
      -- 
    ca_5267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2055_inst_ack_1, ack => convTransposeB_CP_4693_elements(61)); -- 
    rr_5275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(61), ack => type_cast_2065_inst_req_0); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2065_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2065_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2065_Sample/ra
      -- 
    ra_5276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2065_inst_ack_0, ack => convTransposeB_CP_4693_elements(62)); -- 
    -- CP-element group 63:  branch  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (13) 
      -- CP-element group 63: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071__exit__
      -- CP-element group 63: 	 branch_block_stmt_1762/if_stmt_2072__entry__
      -- CP-element group 63: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/$exit
      -- CP-element group 63: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2065_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2065_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_1762/assign_stmt_2036_to_assign_stmt_2071/type_cast_2065_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_1762/if_stmt_2072_dead_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1762/if_stmt_2072_eval_test/$entry
      -- CP-element group 63: 	 branch_block_stmt_1762/if_stmt_2072_eval_test/$exit
      -- CP-element group 63: 	 branch_block_stmt_1762/if_stmt_2072_eval_test/branch_req
      -- CP-element group 63: 	 branch_block_stmt_1762/R_cmp132_2073_place
      -- CP-element group 63: 	 branch_block_stmt_1762/if_stmt_2072_if_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1762/if_stmt_2072_else_link/$entry
      -- 
    ca_5281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2065_inst_ack_1, ack => convTransposeB_CP_4693_elements(63)); -- 
    branch_req_5289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(63), ack => if_stmt_2072_branch_req_0); -- 
    -- CP-element group 64:  merge  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (15) 
      -- CP-element group 64: 	 branch_block_stmt_1762/merge_stmt_2078__exit__
      -- CP-element group 64: 	 branch_block_stmt_1762/assign_stmt_2083__entry__
      -- CP-element group 64: 	 branch_block_stmt_1762/if_stmt_2072_if_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_1762/if_stmt_2072_if_link/if_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_1762/ifx_xelse_whilex_xend
      -- CP-element group 64: 	 branch_block_stmt_1762/assign_stmt_2083/$entry
      -- CP-element group 64: 	 branch_block_stmt_1762/assign_stmt_2083/WPIPE_Block1_done_2080_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_1762/assign_stmt_2083/WPIPE_Block1_done_2080_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1762/assign_stmt_2083/WPIPE_Block1_done_2080_Sample/req
      -- CP-element group 64: 	 branch_block_stmt_1762/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_1762/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 64: 	 branch_block_stmt_1762/merge_stmt_2078_PhiReqMerge
      -- CP-element group 64: 	 branch_block_stmt_1762/merge_stmt_2078_PhiAck/$entry
      -- CP-element group 64: 	 branch_block_stmt_1762/merge_stmt_2078_PhiAck/$exit
      -- CP-element group 64: 	 branch_block_stmt_1762/merge_stmt_2078_PhiAck/dummy
      -- 
    if_choice_transition_5294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2072_branch_ack_1, ack => convTransposeB_CP_4693_elements(64)); -- 
    req_5311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(64), ack => WPIPE_Block1_done_2080_inst_req_0); -- 
    -- CP-element group 65:  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	73 
    -- CP-element group 65: 	74 
    -- CP-element group 65: 	76 
    -- CP-element group 65: 	77 
    -- CP-element group 65:  members (20) 
      -- CP-element group 65: 	 branch_block_stmt_1762/if_stmt_2072_else_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_1762/if_stmt_2072_else_link/else_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 65: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/$entry
      -- CP-element group 65: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1853/$entry
      -- CP-element group 65: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1853/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1853/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1853/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1853/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1853/SplitProtocol/Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/$entry
      -- CP-element group 65: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1860/$entry
      -- CP-element group 65: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1860/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1860/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1860/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1860/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1860/SplitProtocol/Update/cr
      -- 
    else_choice_transition_5298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2072_branch_ack_0, ack => convTransposeB_CP_4693_elements(65)); -- 
    rr_5370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(65), ack => type_cast_1853_inst_req_0); -- 
    cr_5375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(65), ack => type_cast_1853_inst_req_1); -- 
    rr_5393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(65), ack => type_cast_1860_inst_req_0); -- 
    cr_5398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(65), ack => type_cast_1860_inst_req_1); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_1762/assign_stmt_2083/WPIPE_Block1_done_2080_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1762/assign_stmt_2083/WPIPE_Block1_done_2080_update_start_
      -- CP-element group 66: 	 branch_block_stmt_1762/assign_stmt_2083/WPIPE_Block1_done_2080_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1762/assign_stmt_2083/WPIPE_Block1_done_2080_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_1762/assign_stmt_2083/WPIPE_Block1_done_2080_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1762/assign_stmt_2083/WPIPE_Block1_done_2080_Update/req
      -- 
    ack_5312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2080_inst_ack_0, ack => convTransposeB_CP_4693_elements(66)); -- 
    req_5316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(66), ack => WPIPE_Block1_done_2080_inst_req_1); -- 
    -- CP-element group 67:  transition  place  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (16) 
      -- CP-element group 67: 	 $exit
      -- CP-element group 67: 	 branch_block_stmt_1762/branch_block_stmt_1762__exit__
      -- CP-element group 67: 	 branch_block_stmt_1762/$exit
      -- CP-element group 67: 	 branch_block_stmt_1762/assign_stmt_2083__exit__
      -- CP-element group 67: 	 branch_block_stmt_1762/return__
      -- CP-element group 67: 	 branch_block_stmt_1762/merge_stmt_2085__exit__
      -- CP-element group 67: 	 branch_block_stmt_1762/assign_stmt_2083/$exit
      -- CP-element group 67: 	 branch_block_stmt_1762/assign_stmt_2083/WPIPE_Block1_done_2080_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1762/assign_stmt_2083/WPIPE_Block1_done_2080_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1762/assign_stmt_2083/WPIPE_Block1_done_2080_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_1762/return___PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_1762/return___PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_1762/merge_stmt_2085_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_1762/merge_stmt_2085_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_1762/merge_stmt_2085_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_1762/merge_stmt_2085_PhiAck/dummy
      -- 
    ack_5317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2080_inst_ack_1, ack => convTransposeB_CP_4693_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	31 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1851/SplitProtocol/Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1851/SplitProtocol/Sample/ra
      -- 
    ra_5337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1851_inst_ack_0, ack => convTransposeB_CP_4693_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	31 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1851/SplitProtocol/Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1851/SplitProtocol/Update/ca
      -- 
    ca_5342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1851_inst_ack_1, ack => convTransposeB_CP_4693_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (5) 
      -- CP-element group 70: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/$exit
      -- CP-element group 70: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/$exit
      -- CP-element group 70: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1851/$exit
      -- CP-element group 70: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1851/SplitProtocol/$exit
      -- CP-element group 70: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_req
      -- 
    phi_stmt_1848_req_5343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1848_req_5343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(70), ack => phi_stmt_1848_req_0); -- 
    convTransposeB_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4693_elements(68) & convTransposeB_CP_4693_elements(69);
      gj_convTransposeB_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4693_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  transition  output  delay-element  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	31 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/$exit
      -- CP-element group 71: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/$exit
      -- CP-element group 71: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1858_konst_delay_trans
      -- CP-element group 71: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/phi_stmt_1854_req
      -- 
    phi_stmt_1854_req_5351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1854_req_5351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(71), ack => phi_stmt_1854_req_0); -- 
    -- Element group convTransposeB_CP_4693_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => convTransposeB_CP_4693_elements(31), ack => convTransposeB_CP_4693_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  join  transition  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	80 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1762/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4693_elements(70) & convTransposeB_CP_4693_elements(71);
      gj_convTransposeB_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4693_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	65 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1853/SplitProtocol/Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1853/SplitProtocol/Sample/ra
      -- 
    ra_5371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1853_inst_ack_0, ack => convTransposeB_CP_4693_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	65 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1853/SplitProtocol/Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1853/SplitProtocol/Update/ca
      -- 
    ca_5376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1853_inst_ack_1, ack => convTransposeB_CP_4693_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	79 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/$exit
      -- CP-element group 75: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/$exit
      -- CP-element group 75: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1853/$exit
      -- CP-element group 75: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_sources/type_cast_1853/SplitProtocol/$exit
      -- CP-element group 75: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1848/phi_stmt_1848_req
      -- 
    phi_stmt_1848_req_5377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1848_req_5377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(75), ack => phi_stmt_1848_req_1); -- 
    convTransposeB_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4693_elements(73) & convTransposeB_CP_4693_elements(74);
      gj_convTransposeB_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4693_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	65 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1860/SplitProtocol/Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1860/SplitProtocol/Sample/ra
      -- 
    ra_5394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1860_inst_ack_0, ack => convTransposeB_CP_4693_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	65 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1860/SplitProtocol/Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1860/SplitProtocol/Update/ca
      -- 
    ca_5399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1860_inst_ack_1, ack => convTransposeB_CP_4693_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/$exit
      -- CP-element group 78: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/$exit
      -- CP-element group 78: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1860/$exit
      -- CP-element group 78: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1860/SplitProtocol/$exit
      -- CP-element group 78: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1854/phi_stmt_1854_req
      -- 
    phi_stmt_1854_req_5400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1854_req_5400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(78), ack => phi_stmt_1854_req_1); -- 
    convTransposeB_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4693_elements(76) & convTransposeB_CP_4693_elements(77);
      gj_convTransposeB_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4693_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	75 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1762/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4693_elements(75) & convTransposeB_CP_4693_elements(78);
      gj_convTransposeB_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4693_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  merge  fork  transition  place  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	72 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1762/merge_stmt_1847_PhiReqMerge
      -- CP-element group 80: 	 branch_block_stmt_1762/merge_stmt_1847_PhiAck/$entry
      -- 
    convTransposeB_CP_4693_elements(80) <= OrReduce(convTransposeB_CP_4693_elements(72) & convTransposeB_CP_4693_elements(79));
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_1762/merge_stmt_1847_PhiAck/phi_stmt_1848_ack
      -- 
    phi_stmt_1848_ack_5405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1848_ack_0, ack => convTransposeB_CP_4693_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_1762/merge_stmt_1847_PhiAck/phi_stmt_1854_ack
      -- 
    phi_stmt_1854_ack_5406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1854_ack_0, ack => convTransposeB_CP_4693_elements(82)); -- 
    -- CP-element group 83:  join  transition  place  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	87 
    -- CP-element group 83:  members (10) 
      -- CP-element group 83: 	 branch_block_stmt_1762/merge_stmt_1847__exit__
      -- CP-element group 83: 	 branch_block_stmt_1762/assign_stmt_1866_to_assign_stmt_1911__entry__
      -- CP-element group 83: 	 branch_block_stmt_1762/assign_stmt_1866_to_assign_stmt_1911__exit__
      -- CP-element group 83: 	 branch_block_stmt_1762/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 83: 	 branch_block_stmt_1762/assign_stmt_1866_to_assign_stmt_1911/$entry
      -- CP-element group 83: 	 branch_block_stmt_1762/assign_stmt_1866_to_assign_stmt_1911/$exit
      -- CP-element group 83: 	 branch_block_stmt_1762/merge_stmt_1847_PhiAck/$exit
      -- CP-element group 83: 	 branch_block_stmt_1762/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 83: 	 branch_block_stmt_1762/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1914/$entry
      -- CP-element group 83: 	 branch_block_stmt_1762/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/$entry
      -- 
    convTransposeB_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4693_elements(81) & convTransposeB_CP_4693_elements(82);
      gj_convTransposeB_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4693_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	56 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/type_cast_1917/SplitProtocol/Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_1762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/type_cast_1917/SplitProtocol/Sample/ra
      -- 
    ra_5426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1917_inst_ack_0, ack => convTransposeB_CP_4693_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	56 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/type_cast_1917/SplitProtocol/Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_1762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/type_cast_1917/SplitProtocol/Update/ca
      -- 
    ca_5431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1917_inst_ack_1, ack => convTransposeB_CP_4693_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_1762/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 86: 	 branch_block_stmt_1762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1914/$exit
      -- CP-element group 86: 	 branch_block_stmt_1762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_1762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/type_cast_1917/$exit
      -- CP-element group 86: 	 branch_block_stmt_1762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/type_cast_1917/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_1762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1914/phi_stmt_1914_req
      -- 
    phi_stmt_1914_req_5432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1914_req_5432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(86), ack => phi_stmt_1914_req_0); -- 
    convTransposeB_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4693_elements(84) & convTransposeB_CP_4693_elements(85);
      gj_convTransposeB_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4693_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  output  delay-element  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	83 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_1762/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 87: 	 branch_block_stmt_1762/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1914/$exit
      -- CP-element group 87: 	 branch_block_stmt_1762/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/$exit
      -- CP-element group 87: 	 branch_block_stmt_1762/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/type_cast_1920_konst_delay_trans
      -- CP-element group 87: 	 branch_block_stmt_1762/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1914/phi_stmt_1914_req
      -- 
    phi_stmt_1914_req_5443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1914_req_5443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(87), ack => phi_stmt_1914_req_1); -- 
    -- Element group convTransposeB_CP_4693_elements(87) is a control-delay.
    cp_element_87_delay: control_delay_element  generic map(name => " 87_delay", delay_value => 1)  port map(req => convTransposeB_CP_4693_elements(83), ack => convTransposeB_CP_4693_elements(87), clk => clk, reset =>reset);
    -- CP-element group 88:  merge  transition  place  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1762/merge_stmt_1913_PhiReqMerge
      -- CP-element group 88: 	 branch_block_stmt_1762/merge_stmt_1913_PhiAck/$entry
      -- 
    convTransposeB_CP_4693_elements(88) <= OrReduce(convTransposeB_CP_4693_elements(86) & convTransposeB_CP_4693_elements(87));
    -- CP-element group 89:  fork  transition  place  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	32 
    -- CP-element group 89: 	33 
    -- CP-element group 89: 	35 
    -- CP-element group 89: 	37 
    -- CP-element group 89: 	39 
    -- CP-element group 89: 	41 
    -- CP-element group 89: 	42 
    -- CP-element group 89: 	43 
    -- CP-element group 89: 	45 
    -- CP-element group 89: 	52 
    -- CP-element group 89: 	53 
    -- CP-element group 89: 	54 
    -- CP-element group 89: 	47 
    -- CP-element group 89: 	49 
    -- CP-element group 89:  members (51) 
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015__entry__
      -- CP-element group 89: 	 branch_block_stmt_1762/merge_stmt_1913__exit__
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/$entry
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_final_index_sum_regn_Update/req
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_final_index_sum_regn_update_start
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1962_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1955_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1961_final_index_sum_regn_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1955_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1941_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1941_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1962_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1962_complete/req
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1941_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1941_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1941_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1955_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1941_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_Update/word_access_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_Update/word_access_complete/word_0/$entry
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1966_Update/word_access_complete/word_0/cr
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1971_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1971_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1971_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1971_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1971_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1971_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1985_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1985_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_1985_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1992_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_final_index_sum_regn_update_start
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_final_index_sum_regn_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/array_obj_ref_1991_final_index_sum_regn_Update/req
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1992_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/addr_of_1992_complete/req
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_Update/word_access_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_Update/word_access_complete/word_0/$entry
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/ptr_deref_1995_Update/word_access_complete/word_0/cr
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_2001_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_2001_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_2001_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_2001_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_2001_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1762/assign_stmt_1927_to_assign_stmt_2015/type_cast_2001_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1762/merge_stmt_1913_PhiAck/$exit
      -- CP-element group 89: 	 branch_block_stmt_1762/merge_stmt_1913_PhiAck/phi_stmt_1914_ack
      -- 
    phi_stmt_1914_ack_5448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1914_ack_0, ack => convTransposeB_CP_4693_elements(89)); -- 
    req_5010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(89), ack => array_obj_ref_1961_index_offset_req_1); -- 
    cr_4979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(89), ack => type_cast_1955_inst_req_1); -- 
    cr_4965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(89), ack => type_cast_1941_inst_req_1); -- 
    req_5025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(89), ack => addr_of_1962_final_reg_req_1); -- 
    rr_4960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(89), ack => type_cast_1941_inst_req_0); -- 
    cr_5070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(89), ack => ptr_deref_1966_load_0_req_1); -- 
    rr_5084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(89), ack => type_cast_1971_inst_req_0); -- 
    cr_5089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(89), ack => type_cast_1971_inst_req_1); -- 
    cr_5103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(89), ack => type_cast_1985_inst_req_1); -- 
    req_5134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(89), ack => array_obj_ref_1991_index_offset_req_1); -- 
    req_5149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(89), ack => addr_of_1992_final_reg_req_1); -- 
    cr_5199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(89), ack => ptr_deref_1995_store_0_req_1); -- 
    rr_5208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(89), ack => type_cast_2001_inst_req_0); -- 
    cr_5213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4693_elements(89), ack => type_cast_2001_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1949_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1979_wire : std_logic_vector(31 downto 0);
    signal R_idxprom96_1990_resized : std_logic_vector(13 downto 0);
    signal R_idxprom96_1990_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1960_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1960_scaled : std_logic_vector(13 downto 0);
    signal add101_2008 : std_logic_vector(31 downto 0);
    signal add43_1932 : std_logic_vector(15 downto 0);
    signal add87_1937 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1961_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1961_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1961_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1961_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1961_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1961_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1991_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1991_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1991_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1991_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1991_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1991_root_address : std_logic_vector(13 downto 0);
    signal arrayidx91_1963 : std_logic_vector(31 downto 0);
    signal arrayidx97_1993 : std_logic_vector(31 downto 0);
    signal call11_1783 : std_logic_vector(15 downto 0);
    signal call13_1786 : std_logic_vector(15 downto 0);
    signal call14_1789 : std_logic_vector(15 downto 0);
    signal call15_1792 : std_logic_vector(15 downto 0);
    signal call17_1795 : std_logic_vector(15 downto 0);
    signal call19_1798 : std_logic_vector(15 downto 0);
    signal call1_1768 : std_logic_vector(15 downto 0);
    signal call3_1771 : std_logic_vector(15 downto 0);
    signal call5_1774 : std_logic_vector(15 downto 0);
    signal call7_1777 : std_logic_vector(15 downto 0);
    signal call9_1780 : std_logic_vector(15 downto 0);
    signal call_1765 : std_logic_vector(15 downto 0);
    signal cmp116_2046 : std_logic_vector(0 downto 0);
    signal cmp132_2071 : std_logic_vector(0 downto 0);
    signal cmp_2015 : std_logic_vector(0 downto 0);
    signal conv100_2002 : std_logic_vector(31 downto 0);
    signal conv104_1809 : std_logic_vector(31 downto 0);
    signal conv112_2041 : std_logic_vector(31 downto 0);
    signal conv115_1813 : std_logic_vector(31 downto 0);
    signal conv127_2066 : std_logic_vector(31 downto 0);
    signal conv130_1817 : std_logic_vector(31 downto 0);
    signal conv90_1942 : std_logic_vector(31 downto 0);
    signal conv94_1972 : std_logic_vector(31 downto 0);
    signal div131_1823 : std_logic_vector(31 downto 0);
    signal div_1805 : std_logic_vector(15 downto 0);
    signal idxprom96_1986 : std_logic_vector(63 downto 0);
    signal idxprom_1956 : std_logic_vector(63 downto 0);
    signal inc120_2056 : std_logic_vector(15 downto 0);
    signal inc_2036 : std_logic_vector(15 downto 0);
    signal indvar_1914 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2028 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_2061 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_1854 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_1848 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2052 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1927 : std_logic_vector(15 downto 0);
    signal ptr_deref_1966_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1966_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1966_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1966_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1966_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1995_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1995_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1995_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1995_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1995_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1995_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr95_1981 : std_logic_vector(31 downto 0);
    signal shr_1951 : std_logic_vector(31 downto 0);
    signal tmp10_1911 : std_logic_vector(15 downto 0);
    signal tmp159_1866 : std_logic_vector(15 downto 0);
    signal tmp160_1871 : std_logic_vector(15 downto 0);
    signal tmp161_1876 : std_logic_vector(15 downto 0);
    signal tmp1_1834 : std_logic_vector(15 downto 0);
    signal tmp2_1881 : std_logic_vector(15 downto 0);
    signal tmp3_1886 : std_logic_vector(15 downto 0);
    signal tmp4_1840 : std_logic_vector(15 downto 0);
    signal tmp5_1845 : std_logic_vector(15 downto 0);
    signal tmp6_1891 : std_logic_vector(15 downto 0);
    signal tmp7_1896 : std_logic_vector(15 downto 0);
    signal tmp8_1901 : std_logic_vector(15 downto 0);
    signal tmp92_1967 : std_logic_vector(63 downto 0);
    signal tmp9_1906 : std_logic_vector(15 downto 0);
    signal tmp_1829 : std_logic_vector(15 downto 0);
    signal type_cast_1803_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1821_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1827_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1838_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1851_wire : std_logic_vector(15 downto 0);
    signal type_cast_1853_wire : std_logic_vector(15 downto 0);
    signal type_cast_1858_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1860_wire : std_logic_vector(15 downto 0);
    signal type_cast_1917_wire : std_logic_vector(15 downto 0);
    signal type_cast_1920_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1925_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1940_wire : std_logic_vector(31 downto 0);
    signal type_cast_1945_wire : std_logic_vector(31 downto 0);
    signal type_cast_1948_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1954_wire : std_logic_vector(63 downto 0);
    signal type_cast_1970_wire : std_logic_vector(31 downto 0);
    signal type_cast_1975_wire : std_logic_vector(31 downto 0);
    signal type_cast_1978_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1984_wire : std_logic_vector(63 downto 0);
    signal type_cast_2000_wire : std_logic_vector(31 downto 0);
    signal type_cast_2006_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2011_wire : std_logic_vector(31 downto 0);
    signal type_cast_2013_wire : std_logic_vector(31 downto 0);
    signal type_cast_2026_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2034_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2039_wire : std_logic_vector(31 downto 0);
    signal type_cast_2064_wire : std_logic_vector(31 downto 0);
    signal type_cast_2082_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_1961_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1961_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1961_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1961_resized_base_address <= "00000000000000";
    array_obj_ref_1991_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1991_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1991_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1991_resized_base_address <= "00000000000000";
    ptr_deref_1966_word_offset_0 <= "00000000000000";
    ptr_deref_1995_word_offset_0 <= "00000000000000";
    type_cast_1803_wire_constant <= "0000000000000001";
    type_cast_1821_wire_constant <= "00000000000000000000000000000001";
    type_cast_1827_wire_constant <= "1111111111111111";
    type_cast_1838_wire_constant <= "1111111111111111";
    type_cast_1858_wire_constant <= "0000000000000000";
    type_cast_1920_wire_constant <= "0000000000000000";
    type_cast_1925_wire_constant <= "0000000000000100";
    type_cast_1948_wire_constant <= "00000000000000000000000000000010";
    type_cast_1978_wire_constant <= "00000000000000000000000000000010";
    type_cast_2006_wire_constant <= "00000000000000000000000000000100";
    type_cast_2026_wire_constant <= "0000000000000001";
    type_cast_2034_wire_constant <= "0000000000000001";
    type_cast_2082_wire_constant <= "0000000000000001";
    phi_stmt_1848: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1851_wire & type_cast_1853_wire;
      req <= phi_stmt_1848_req_0 & phi_stmt_1848_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1848",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1848_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_1848,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1848
    phi_stmt_1854: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1858_wire_constant & type_cast_1860_wire;
      req <= phi_stmt_1854_req_0 & phi_stmt_1854_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1854",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1854_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_1854,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1854
    phi_stmt_1914: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1917_wire & type_cast_1920_wire_constant;
      req <= phi_stmt_1914_req_0 & phi_stmt_1914_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1914",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1914_ack_0,
          idata => idata,
          odata => indvar_1914,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1914
    -- flow-through select operator MUX_2051_inst
    input_dim1x_x2_2052 <= div_1805 when (cmp116_2046(0) /=  '0') else inc_2036;
    addr_of_1962_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1962_final_reg_req_0;
      addr_of_1962_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1962_final_reg_req_1;
      addr_of_1962_final_reg_ack_1<= rack(0);
      addr_of_1962_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1962_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1961_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx91_1963,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1992_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1992_final_reg_req_0;
      addr_of_1992_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1992_final_reg_req_1;
      addr_of_1992_final_reg_ack_1<= rack(0);
      addr_of_1992_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1992_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1991_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx97_1993,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1808_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1808_inst_req_0;
      type_cast_1808_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1808_inst_req_1;
      type_cast_1808_inst_ack_1<= rack(0);
      type_cast_1808_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1808_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1771,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_1809,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1812_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1812_inst_req_0;
      type_cast_1812_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1812_inst_req_1;
      type_cast_1812_inst_ack_1<= rack(0);
      type_cast_1812_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1812_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_1768,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_1813,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1816_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1816_inst_req_0;
      type_cast_1816_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1816_inst_req_1;
      type_cast_1816_inst_ack_1<= rack(0);
      type_cast_1816_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1816_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1765,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv130_1817,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1851_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1851_inst_req_0;
      type_cast_1851_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1851_inst_req_1;
      type_cast_1851_inst_ack_1<= rack(0);
      type_cast_1851_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1851_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_1805,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1851_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1853_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1853_inst_req_0;
      type_cast_1853_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1853_inst_req_1;
      type_cast_1853_inst_ack_1<= rack(0);
      type_cast_1853_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1853_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2052,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1853_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1860_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1860_inst_req_0;
      type_cast_1860_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1860_inst_req_1;
      type_cast_1860_inst_ack_1<= rack(0);
      type_cast_1860_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1860_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_2061,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1860_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1917_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1917_inst_req_0;
      type_cast_1917_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1917_inst_req_1;
      type_cast_1917_inst_ack_1<= rack(0);
      type_cast_1917_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1917_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2028,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1917_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1941_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1941_inst_req_0;
      type_cast_1941_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1941_inst_req_1;
      type_cast_1941_inst_ack_1<= rack(0);
      type_cast_1941_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1941_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1940_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_1942,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1945_inst
    process(conv90_1942) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv90_1942(31 downto 0);
      type_cast_1945_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1950_inst
    process(ASHR_i32_i32_1949_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1949_wire(31 downto 0);
      shr_1951 <= tmp_var; -- 
    end process;
    type_cast_1955_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1955_inst_req_0;
      type_cast_1955_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1955_inst_req_1;
      type_cast_1955_inst_ack_1<= rack(0);
      type_cast_1955_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1955_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1954_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1956,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1971_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1971_inst_req_0;
      type_cast_1971_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1971_inst_req_1;
      type_cast_1971_inst_ack_1<= rack(0);
      type_cast_1971_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1971_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1970_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_1972,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1975_inst
    process(conv94_1972) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv94_1972(31 downto 0);
      type_cast_1975_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1980_inst
    process(ASHR_i32_i32_1979_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1979_wire(31 downto 0);
      shr95_1981 <= tmp_var; -- 
    end process;
    type_cast_1985_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1985_inst_req_0;
      type_cast_1985_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1985_inst_req_1;
      type_cast_1985_inst_ack_1<= rack(0);
      type_cast_1985_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1985_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1984_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom96_1986,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2001_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2001_inst_req_0;
      type_cast_2001_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2001_inst_req_1;
      type_cast_2001_inst_ack_1<= rack(0);
      type_cast_2001_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2001_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2000_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv100_2002,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2011_inst
    process(add101_2008) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add101_2008(31 downto 0);
      type_cast_2011_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2013_inst
    process(conv104_1809) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv104_1809(31 downto 0);
      type_cast_2013_wire <= tmp_var; -- 
    end process;
    type_cast_2040_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2040_inst_req_0;
      type_cast_2040_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2040_inst_req_1;
      type_cast_2040_inst_ack_1<= rack(0);
      type_cast_2040_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2040_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2039_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_2041,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2055_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2055_inst_req_0;
      type_cast_2055_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2055_inst_req_1;
      type_cast_2055_inst_ack_1<= rack(0);
      type_cast_2055_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2055_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp116_2046,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc120_2056,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2065_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2065_inst_req_0;
      type_cast_2065_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2065_inst_req_1;
      type_cast_2065_inst_ack_1<= rack(0);
      type_cast_2065_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2065_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2064_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv127_2066,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1961_index_1_rename
    process(R_idxprom_1960_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1960_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1960_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1961_index_1_resize
    process(idxprom_1956) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1956;
      ov := iv(13 downto 0);
      R_idxprom_1960_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1961_root_address_inst
    process(array_obj_ref_1961_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1961_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1961_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1991_index_1_rename
    process(R_idxprom96_1990_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom96_1990_resized;
      ov(13 downto 0) := iv;
      R_idxprom96_1990_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1991_index_1_resize
    process(idxprom96_1986) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom96_1986;
      ov := iv(13 downto 0);
      R_idxprom96_1990_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1991_root_address_inst
    process(array_obj_ref_1991_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1991_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1991_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1966_addr_0
    process(ptr_deref_1966_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1966_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1966_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1966_base_resize
    process(arrayidx91_1963) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx91_1963;
      ov := iv(13 downto 0);
      ptr_deref_1966_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1966_gather_scatter
    process(ptr_deref_1966_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1966_data_0;
      ov(63 downto 0) := iv;
      tmp92_1967 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1966_root_address_inst
    process(ptr_deref_1966_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1966_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1966_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1995_addr_0
    process(ptr_deref_1995_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1995_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1995_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1995_base_resize
    process(arrayidx97_1993) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx97_1993;
      ov := iv(13 downto 0);
      ptr_deref_1995_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1995_gather_scatter
    process(tmp92_1967) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp92_1967;
      ov(63 downto 0) := iv;
      ptr_deref_1995_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1995_root_address_inst
    process(ptr_deref_1995_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1995_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1995_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2016_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2015;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2016_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2016_branch_req_0,
          ack0 => if_stmt_2016_branch_ack_0,
          ack1 => if_stmt_2016_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2072_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp132_2071;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2072_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2072_branch_req_0,
          ack0 => if_stmt_2072_branch_ack_0,
          ack1 => if_stmt_2072_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1828_inst
    process(call9_1780) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1780, type_cast_1827_wire_constant, tmp_var);
      tmp_1829 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1839_inst
    process(call7_1777) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1777, type_cast_1838_wire_constant, tmp_var);
      tmp4_1840 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1870_inst
    process(input_dim1x_x1x_xph_1848, tmp159_1866) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1848, tmp159_1866, tmp_var);
      tmp160_1871 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1885_inst
    process(tmp1_1834, tmp2_1881) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp1_1834, tmp2_1881, tmp_var);
      tmp3_1886 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1895_inst
    process(tmp5_1845, tmp6_1891) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp5_1845, tmp6_1891, tmp_var);
      tmp7_1896 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1905_inst
    process(tmp3_1886, tmp8_1901) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_1886, tmp8_1901, tmp_var);
      tmp9_1906 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1931_inst
    process(tmp161_1876, input_dim2x_x1_1927) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp161_1876, input_dim2x_x1_1927, tmp_var);
      add43_1932 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1936_inst
    process(tmp10_1911, input_dim2x_x1_1927) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp10_1911, input_dim2x_x1_1927, tmp_var);
      add87_1937 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2027_inst
    process(indvar_1914) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1914, type_cast_2026_wire_constant, tmp_var);
      indvarx_xnext_2028 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2035_inst
    process(input_dim1x_x1x_xph_1848) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1848, type_cast_2034_wire_constant, tmp_var);
      inc_2036 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2060_inst
    process(inc120_2056, input_dim0x_x2x_xph_1854) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc120_2056, input_dim0x_x2x_xph_1854, tmp_var);
      input_dim0x_x0_2061 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2007_inst
    process(conv100_2002) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv100_2002, type_cast_2006_wire_constant, tmp_var);
      add101_2008 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1949_inst
    process(type_cast_1945_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1945_wire, type_cast_1948_wire_constant, tmp_var);
      ASHR_i32_i32_1949_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1979_inst
    process(type_cast_1975_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1975_wire, type_cast_1978_wire_constant, tmp_var);
      ASHR_i32_i32_1979_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2045_inst
    process(conv112_2041, conv115_1813) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv112_2041, conv115_1813, tmp_var);
      cmp116_2046 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2070_inst
    process(conv127_2066, div131_1823) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv127_2066, div131_1823, tmp_var);
      cmp132_2071 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1804_inst
    process(call1_1768) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call1_1768, type_cast_1803_wire_constant, tmp_var);
      div_1805 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1822_inst
    process(conv130_1817) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv130_1817, type_cast_1821_wire_constant, tmp_var);
      div131_1823 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1865_inst
    process(call1_1768, input_dim0x_x2x_xph_1854) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call1_1768, input_dim0x_x2x_xph_1854, tmp_var);
      tmp159_1866 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1875_inst
    process(call3_1771, tmp160_1871) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call3_1771, tmp160_1871, tmp_var);
      tmp161_1876 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1880_inst
    process(call13_1786, input_dim1x_x1x_xph_1848) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_1786, input_dim1x_x1x_xph_1848, tmp_var);
      tmp2_1881 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1890_inst
    process(call13_1786, input_dim0x_x2x_xph_1854) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_1786, input_dim0x_x2x_xph_1854, tmp_var);
      tmp6_1891 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1900_inst
    process(call17_1795, tmp7_1896) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call17_1795, tmp7_1896, tmp_var);
      tmp8_1901 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1910_inst
    process(call19_1798, tmp9_1906) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call19_1798, tmp9_1906, tmp_var);
      tmp10_1911 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1926_inst
    process(indvar_1914) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1914, type_cast_1925_wire_constant, tmp_var);
      input_dim2x_x1_1927 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2014_inst
    process(type_cast_2011_wire, type_cast_2013_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2011_wire, type_cast_2013_wire, tmp_var);
      cmp_2015 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1833_inst
    process(tmp_1829, call14_1789) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp_1829, call14_1789, tmp_var);
      tmp1_1834 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1844_inst
    process(tmp4_1840, call14_1789) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp4_1840, call14_1789, tmp_var);
      tmp5_1845 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_1961_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1960_scaled;
      array_obj_ref_1961_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1961_index_offset_req_0;
      array_obj_ref_1961_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1961_index_offset_req_1;
      array_obj_ref_1961_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_1991_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom96_1990_scaled;
      array_obj_ref_1991_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1991_index_offset_req_0;
      array_obj_ref_1991_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1991_index_offset_req_1;
      array_obj_ref_1991_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- unary operator type_cast_1940_inst
    process(add43_1932) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add43_1932, tmp_var);
      type_cast_1940_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1954_inst
    process(shr_1951) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1951, tmp_var);
      type_cast_1954_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1970_inst
    process(add87_1937) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add87_1937, tmp_var);
      type_cast_1970_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1984_inst
    process(shr95_1981) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr95_1981, tmp_var);
      type_cast_1984_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2000_inst
    process(input_dim2x_x1_1927) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_1927, tmp_var);
      type_cast_2000_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2039_inst
    process(inc_2036) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2036, tmp_var);
      type_cast_2039_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2064_inst
    process(input_dim0x_x0_2061) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x0_2061, tmp_var);
      type_cast_2064_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1966_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1966_load_0_req_0;
      ptr_deref_1966_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1966_load_0_req_1;
      ptr_deref_1966_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1966_word_address_0;
      ptr_deref_1966_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1995_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1995_store_0_req_0;
      ptr_deref_1995_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1995_store_0_req_1;
      ptr_deref_1995_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1995_word_address_0;
      data_in <= ptr_deref_1995_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1797_inst RPIPE_Block1_start_1794_inst RPIPE_Block1_start_1791_inst RPIPE_Block1_start_1788_inst RPIPE_Block1_start_1785_inst RPIPE_Block1_start_1782_inst RPIPE_Block1_start_1779_inst RPIPE_Block1_start_1776_inst RPIPE_Block1_start_1773_inst RPIPE_Block1_start_1770_inst RPIPE_Block1_start_1767_inst RPIPE_Block1_start_1764_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(191 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 11 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 11 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant outBUFs : IntegerArray(11 downto 0) := (11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      reqL_unguarded(11) <= RPIPE_Block1_start_1797_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block1_start_1794_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block1_start_1791_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block1_start_1788_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block1_start_1785_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block1_start_1782_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block1_start_1779_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block1_start_1776_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block1_start_1773_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block1_start_1770_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block1_start_1767_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block1_start_1764_inst_req_0;
      RPIPE_Block1_start_1797_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block1_start_1794_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block1_start_1791_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block1_start_1788_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block1_start_1785_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block1_start_1782_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block1_start_1779_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block1_start_1776_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block1_start_1773_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block1_start_1770_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block1_start_1767_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block1_start_1764_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(11) <= RPIPE_Block1_start_1797_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block1_start_1794_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block1_start_1791_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block1_start_1788_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block1_start_1785_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block1_start_1782_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block1_start_1779_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block1_start_1776_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block1_start_1773_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block1_start_1770_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block1_start_1767_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block1_start_1764_inst_req_1;
      RPIPE_Block1_start_1797_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block1_start_1794_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block1_start_1791_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block1_start_1788_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block1_start_1785_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block1_start_1782_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block1_start_1779_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block1_start_1776_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block1_start_1773_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block1_start_1770_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block1_start_1767_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block1_start_1764_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      call19_1798 <= data_out(191 downto 176);
      call17_1795 <= data_out(175 downto 160);
      call15_1792 <= data_out(159 downto 144);
      call14_1789 <= data_out(143 downto 128);
      call13_1786 <= data_out(127 downto 112);
      call11_1783 <= data_out(111 downto 96);
      call9_1780 <= data_out(95 downto 80);
      call7_1777 <= data_out(79 downto 64);
      call5_1774 <= data_out(63 downto 48);
      call3_1771 <= data_out(47 downto 32);
      call1_1768 <= data_out(31 downto 16);
      call_1765 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 12,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_2080_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_2080_inst_req_0;
      WPIPE_Block1_done_2080_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_2080_inst_req_1;
      WPIPE_Block1_done_2080_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2082_wire_constant;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_5489_start: Boolean;
  signal convTransposeC_CP_5489_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_2244_inst_req_1 : boolean;
  signal array_obj_ref_2318_index_offset_ack_1 : boolean;
  signal if_stmt_2400_branch_req_0 : boolean;
  signal type_cast_2393_inst_req_0 : boolean;
  signal WPIPE_Block2_done_2408_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2091_inst_req_0 : boolean;
  signal type_cast_2185_inst_ack_0 : boolean;
  signal type_cast_2187_inst_req_0 : boolean;
  signal phi_stmt_2182_req_0 : boolean;
  signal phi_stmt_2175_req_0 : boolean;
  signal type_cast_2244_inst_ack_1 : boolean;
  signal type_cast_2187_inst_ack_0 : boolean;
  signal if_stmt_2400_branch_ack_1 : boolean;
  signal phi_stmt_2241_req_0 : boolean;
  signal type_cast_2393_inst_ack_0 : boolean;
  signal phi_stmt_2241_ack_0 : boolean;
  signal if_stmt_2343_branch_ack_1 : boolean;
  signal type_cast_2328_inst_req_1 : boolean;
  signal array_obj_ref_2318_index_offset_req_1 : boolean;
  signal if_stmt_2400_branch_ack_0 : boolean;
  signal WPIPE_Block2_done_2408_inst_req_1 : boolean;
  signal if_stmt_2343_branch_req_0 : boolean;
  signal type_cast_2187_inst_req_1 : boolean;
  signal type_cast_2185_inst_req_1 : boolean;
  signal type_cast_2185_inst_ack_1 : boolean;
  signal type_cast_2393_inst_ack_1 : boolean;
  signal WPIPE_Block2_done_2408_inst_req_0 : boolean;
  signal type_cast_2187_inst_ack_1 : boolean;
  signal type_cast_2393_inst_req_1 : boolean;
  signal phi_stmt_2182_req_1 : boolean;
  signal if_stmt_2343_branch_ack_0 : boolean;
  signal array_obj_ref_2318_index_offset_ack_0 : boolean;
  signal type_cast_2376_inst_req_1 : boolean;
  signal type_cast_2376_inst_ack_1 : boolean;
  signal WPIPE_Block2_done_2408_inst_ack_0 : boolean;
  signal type_cast_2328_inst_ack_1 : boolean;
  signal type_cast_2185_inst_req_0 : boolean;
  signal phi_stmt_2241_req_1 : boolean;
  signal RPIPE_Block2_start_2091_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2091_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2091_inst_ack_1 : boolean;
  signal type_cast_2244_inst_ack_0 : boolean;
  signal type_cast_2244_inst_req_0 : boolean;
  signal type_cast_2328_inst_ack_0 : boolean;
  signal type_cast_2328_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2094_inst_req_0 : boolean;
  signal type_cast_2376_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2094_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2094_inst_req_1 : boolean;
  signal type_cast_2376_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2094_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2097_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2097_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2097_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2097_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2100_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2100_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2100_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2100_inst_ack_1 : boolean;
  signal addr_of_2319_final_reg_ack_1 : boolean;
  signal phi_stmt_2182_ack_0 : boolean;
  signal phi_stmt_2175_ack_0 : boolean;
  signal ptr_deref_2322_store_0_ack_1 : boolean;
  signal ptr_deref_2322_store_0_req_1 : boolean;
  signal RPIPE_Block2_start_2103_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2103_inst_ack_0 : boolean;
  signal addr_of_2319_final_reg_req_1 : boolean;
  signal RPIPE_Block2_start_2103_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2103_inst_ack_1 : boolean;
  signal phi_stmt_2175_req_1 : boolean;
  signal type_cast_2181_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2106_inst_req_0 : boolean;
  signal type_cast_2367_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2106_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2106_inst_req_1 : boolean;
  signal type_cast_2367_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2106_inst_ack_1 : boolean;
  signal addr_of_2319_final_reg_ack_0 : boolean;
  signal type_cast_2181_inst_req_1 : boolean;
  signal type_cast_2181_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2109_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2109_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2109_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2109_inst_ack_1 : boolean;
  signal array_obj_ref_2318_index_offset_req_0 : boolean;
  signal type_cast_2181_inst_req_0 : boolean;
  signal ptr_deref_2322_store_0_ack_0 : boolean;
  signal RPIPE_Block2_start_2112_inst_req_0 : boolean;
  signal type_cast_2367_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2112_inst_ack_0 : boolean;
  signal addr_of_2319_final_reg_req_0 : boolean;
  signal RPIPE_Block2_start_2112_inst_req_1 : boolean;
  signal type_cast_2367_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2112_inst_ack_1 : boolean;
  signal ptr_deref_2322_store_0_req_0 : boolean;
  signal RPIPE_Block2_start_2115_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2115_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2115_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2115_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2118_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2118_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2118_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2118_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2121_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2121_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2121_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2121_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2124_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2124_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2124_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2124_inst_ack_1 : boolean;
  signal type_cast_2135_inst_req_0 : boolean;
  signal type_cast_2135_inst_ack_0 : boolean;
  signal type_cast_2135_inst_req_1 : boolean;
  signal type_cast_2135_inst_ack_1 : boolean;
  signal type_cast_2139_inst_req_0 : boolean;
  signal type_cast_2139_inst_ack_0 : boolean;
  signal type_cast_2139_inst_req_1 : boolean;
  signal type_cast_2139_inst_ack_1 : boolean;
  signal type_cast_2149_inst_req_0 : boolean;
  signal type_cast_2149_inst_ack_0 : boolean;
  signal type_cast_2149_inst_req_1 : boolean;
  signal type_cast_2149_inst_ack_1 : boolean;
  signal type_cast_2268_inst_req_0 : boolean;
  signal type_cast_2268_inst_ack_0 : boolean;
  signal type_cast_2268_inst_req_1 : boolean;
  signal type_cast_2268_inst_ack_1 : boolean;
  signal type_cast_2282_inst_req_0 : boolean;
  signal type_cast_2282_inst_ack_0 : boolean;
  signal type_cast_2282_inst_req_1 : boolean;
  signal type_cast_2282_inst_ack_1 : boolean;
  signal array_obj_ref_2288_index_offset_req_0 : boolean;
  signal array_obj_ref_2288_index_offset_ack_0 : boolean;
  signal array_obj_ref_2288_index_offset_req_1 : boolean;
  signal array_obj_ref_2288_index_offset_ack_1 : boolean;
  signal addr_of_2289_final_reg_req_0 : boolean;
  signal addr_of_2289_final_reg_ack_0 : boolean;
  signal addr_of_2289_final_reg_req_1 : boolean;
  signal addr_of_2289_final_reg_ack_1 : boolean;
  signal ptr_deref_2293_load_0_req_0 : boolean;
  signal ptr_deref_2293_load_0_ack_0 : boolean;
  signal ptr_deref_2293_load_0_req_1 : boolean;
  signal ptr_deref_2293_load_0_ack_1 : boolean;
  signal type_cast_2298_inst_req_0 : boolean;
  signal type_cast_2298_inst_ack_0 : boolean;
  signal type_cast_2298_inst_req_1 : boolean;
  signal type_cast_2298_inst_ack_1 : boolean;
  signal type_cast_2312_inst_req_0 : boolean;
  signal type_cast_2312_inst_ack_0 : boolean;
  signal type_cast_2312_inst_req_1 : boolean;
  signal type_cast_2312_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_5489_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5489_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_5489_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5489_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_5489: Block -- control-path 
    signal convTransposeC_CP_5489_elements: BooleanArray(89 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_5489_elements(0) <= convTransposeC_CP_5489_start;
    convTransposeC_CP_5489_symbol <= convTransposeC_CP_5489_elements(67);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2091_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125__entry__
      -- CP-element group 0: 	 branch_block_stmt_2089/$entry
      -- CP-element group 0: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/$entry
      -- CP-element group 0: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2091_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2091_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2089/branch_block_stmt_2089__entry__
      -- CP-element group 0: 	 $entry
      -- 
    rr_5537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(0), ack => RPIPE_Block2_start_2091_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2091_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2091_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2091_update_start_
      -- CP-element group 1: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2091_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2091_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2091_Update/cr
      -- 
    ra_5538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2091_inst_ack_0, ack => convTransposeC_CP_5489_elements(1)); -- 
    cr_5542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(1), ack => RPIPE_Block2_start_2091_inst_req_1); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2091_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2091_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2091_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2094_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2094_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2094_Sample/rr
      -- 
    ca_5543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2091_inst_ack_1, ack => convTransposeC_CP_5489_elements(2)); -- 
    rr_5551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(2), ack => RPIPE_Block2_start_2094_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2094_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2094_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2094_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2094_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2094_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2094_Update/cr
      -- 
    ra_5552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2094_inst_ack_0, ack => convTransposeC_CP_5489_elements(3)); -- 
    cr_5556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(3), ack => RPIPE_Block2_start_2094_inst_req_1); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2094_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2094_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2094_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2097_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2097_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2097_Sample/rr
      -- 
    ca_5557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2094_inst_ack_1, ack => convTransposeC_CP_5489_elements(4)); -- 
    rr_5565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(4), ack => RPIPE_Block2_start_2097_inst_req_0); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2097_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2097_update_start_
      -- CP-element group 5: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2097_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2097_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2097_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2097_Update/cr
      -- 
    ra_5566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2097_inst_ack_0, ack => convTransposeC_CP_5489_elements(5)); -- 
    cr_5570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(5), ack => RPIPE_Block2_start_2097_inst_req_1); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2097_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2097_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2097_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2100_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2100_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2100_Sample/rr
      -- 
    ca_5571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2097_inst_ack_1, ack => convTransposeC_CP_5489_elements(6)); -- 
    rr_5579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(6), ack => RPIPE_Block2_start_2100_inst_req_0); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2100_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2100_update_start_
      -- CP-element group 7: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2100_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2100_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2100_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2100_Update/cr
      -- 
    ra_5580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2100_inst_ack_0, ack => convTransposeC_CP_5489_elements(7)); -- 
    cr_5584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(7), ack => RPIPE_Block2_start_2100_inst_req_1); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2100_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2100_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2100_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2103_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2103_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2103_Sample/rr
      -- 
    ca_5585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2100_inst_ack_1, ack => convTransposeC_CP_5489_elements(8)); -- 
    rr_5593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(8), ack => RPIPE_Block2_start_2103_inst_req_0); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2103_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2103_update_start_
      -- CP-element group 9: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2103_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2103_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2103_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2103_Update/cr
      -- 
    ra_5594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2103_inst_ack_0, ack => convTransposeC_CP_5489_elements(9)); -- 
    cr_5598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(9), ack => RPIPE_Block2_start_2103_inst_req_1); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2103_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2103_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2103_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2106_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2106_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2106_Sample/rr
      -- 
    ca_5599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2103_inst_ack_1, ack => convTransposeC_CP_5489_elements(10)); -- 
    rr_5607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(10), ack => RPIPE_Block2_start_2106_inst_req_0); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2106_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2106_update_start_
      -- CP-element group 11: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2106_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2106_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2106_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2106_Update/cr
      -- 
    ra_5608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2106_inst_ack_0, ack => convTransposeC_CP_5489_elements(11)); -- 
    cr_5612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(11), ack => RPIPE_Block2_start_2106_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2106_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2106_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2106_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2109_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2109_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2109_Sample/rr
      -- 
    ca_5613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2106_inst_ack_1, ack => convTransposeC_CP_5489_elements(12)); -- 
    rr_5621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(12), ack => RPIPE_Block2_start_2109_inst_req_0); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2109_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2109_update_start_
      -- CP-element group 13: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2109_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2109_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2109_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2109_Update/cr
      -- 
    ra_5622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2109_inst_ack_0, ack => convTransposeC_CP_5489_elements(13)); -- 
    cr_5626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(13), ack => RPIPE_Block2_start_2109_inst_req_1); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2109_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2109_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2109_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2112_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2112_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2112_Sample/rr
      -- 
    ca_5627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2109_inst_ack_1, ack => convTransposeC_CP_5489_elements(14)); -- 
    rr_5635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(14), ack => RPIPE_Block2_start_2112_inst_req_0); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2112_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2112_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2112_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2112_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2112_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2112_Update/cr
      -- 
    ra_5636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2112_inst_ack_0, ack => convTransposeC_CP_5489_elements(15)); -- 
    cr_5640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(15), ack => RPIPE_Block2_start_2112_inst_req_1); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2112_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2112_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2112_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2115_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2115_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2115_Sample/rr
      -- 
    ca_5641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2112_inst_ack_1, ack => convTransposeC_CP_5489_elements(16)); -- 
    rr_5649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(16), ack => RPIPE_Block2_start_2115_inst_req_0); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2115_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2115_update_start_
      -- CP-element group 17: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2115_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2115_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2115_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2115_Update/cr
      -- 
    ra_5650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2115_inst_ack_0, ack => convTransposeC_CP_5489_elements(17)); -- 
    cr_5654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(17), ack => RPIPE_Block2_start_2115_inst_req_1); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2115_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2115_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2115_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2118_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2118_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2118_Sample/rr
      -- 
    ca_5655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2115_inst_ack_1, ack => convTransposeC_CP_5489_elements(18)); -- 
    rr_5663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(18), ack => RPIPE_Block2_start_2118_inst_req_0); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2118_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2118_update_start_
      -- CP-element group 19: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2118_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2118_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2118_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2118_Update/cr
      -- 
    ra_5664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2118_inst_ack_0, ack => convTransposeC_CP_5489_elements(19)); -- 
    cr_5668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(19), ack => RPIPE_Block2_start_2118_inst_req_1); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2118_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2118_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2118_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2121_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2121_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2121_Sample/rr
      -- 
    ca_5669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2118_inst_ack_1, ack => convTransposeC_CP_5489_elements(20)); -- 
    rr_5677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(20), ack => RPIPE_Block2_start_2121_inst_req_0); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2121_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2121_update_start_
      -- CP-element group 21: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2121_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2121_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2121_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2121_Update/cr
      -- 
    ra_5678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2121_inst_ack_0, ack => convTransposeC_CP_5489_elements(21)); -- 
    cr_5682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(21), ack => RPIPE_Block2_start_2121_inst_req_1); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2121_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2121_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2121_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2124_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2124_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2124_Sample/rr
      -- 
    ca_5683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2121_inst_ack_1, ack => convTransposeC_CP_5489_elements(22)); -- 
    rr_5691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(22), ack => RPIPE_Block2_start_2124_inst_req_0); -- 
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2124_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2124_update_start_
      -- CP-element group 23: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2124_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2124_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2124_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2124_Update/cr
      -- 
    ra_5692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2124_inst_ack_0, ack => convTransposeC_CP_5489_elements(23)); -- 
    cr_5696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(23), ack => RPIPE_Block2_start_2124_inst_req_1); -- 
    -- CP-element group 24:  fork  transition  place  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	27 
    -- CP-element group 24: 	28 
    -- CP-element group 24: 	29 
    -- CP-element group 24: 	30 
    -- CP-element group 24:  members (25) 
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172__entry__
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125__exit__
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/$exit
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2124_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2124_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2092_to_assign_stmt_2125/RPIPE_Block2_start_2124_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/$entry
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2135_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2135_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2135_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2135_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2135_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2135_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2139_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2139_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2139_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2139_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2139_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2139_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2149_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2149_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2149_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2149_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2149_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2149_Update/cr
      -- 
    ca_5697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2124_inst_ack_1, ack => convTransposeC_CP_5489_elements(24)); -- 
    rr_5708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(24), ack => type_cast_2135_inst_req_0); -- 
    cr_5713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(24), ack => type_cast_2135_inst_req_1); -- 
    rr_5722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(24), ack => type_cast_2139_inst_req_0); -- 
    cr_5727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(24), ack => type_cast_2139_inst_req_1); -- 
    rr_5736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(24), ack => type_cast_2149_inst_req_0); -- 
    cr_5741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(24), ack => type_cast_2149_inst_req_1); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2135_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2135_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2135_Sample/ra
      -- 
    ra_5709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2135_inst_ack_0, ack => convTransposeC_CP_5489_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2135_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2135_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2135_Update/ca
      -- 
    ca_5714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2135_inst_ack_1, ack => convTransposeC_CP_5489_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	24 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2139_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2139_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2139_Sample/ra
      -- 
    ra_5723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2139_inst_ack_0, ack => convTransposeC_CP_5489_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	24 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2139_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2139_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2139_Update/ca
      -- 
    ca_5728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2139_inst_ack_1, ack => convTransposeC_CP_5489_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	24 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2149_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2149_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2149_Sample/ra
      -- 
    ra_5737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2149_inst_ack_0, ack => convTransposeC_CP_5489_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	24 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2149_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2149_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/type_cast_2149_Update/ca
      -- 
    ca_5742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2149_inst_ack_1, ack => convTransposeC_CP_5489_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	68 
    -- CP-element group 31: 	69 
    -- CP-element group 31: 	71 
    -- CP-element group 31:  members (14) 
      -- CP-element group 31: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/$entry
      -- CP-element group 31: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172__exit__
      -- CP-element group 31: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/$entry
      -- CP-element group 31: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/SplitProtocol/Update/cr
      -- CP-element group 31: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/SplitProtocol/Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/$entry
      -- CP-element group 31: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2089/assign_stmt_2132_to_assign_stmt_2172/$exit
      -- 
    cr_6137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(31), ack => type_cast_2185_inst_req_1); -- 
    rr_6132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(31), ack => type_cast_2185_inst_req_0); -- 
    convTransposeC_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5489_elements(26) & convTransposeC_CP_5489_elements(28) & convTransposeC_CP_5489_elements(30);
      gj_convTransposeC_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5489_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	89 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2268_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2268_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2268_Sample/ra
      -- 
    ra_5757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2268_inst_ack_0, ack => convTransposeC_CP_5489_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	89 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2268_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2268_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2268_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2282_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2282_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2282_Sample/rr
      -- 
    ca_5762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2268_inst_ack_1, ack => convTransposeC_CP_5489_elements(33)); -- 
    rr_5770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(33), ack => type_cast_2282_inst_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2282_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2282_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2282_Sample/ra
      -- 
    ra_5771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2282_inst_ack_0, ack => convTransposeC_CP_5489_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	89 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (16) 
      -- CP-element group 35: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2282_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2282_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2282_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_index_resized_1
      -- CP-element group 35: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_index_scaled_1
      -- CP-element group 35: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_index_computed_1
      -- CP-element group 35: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_index_resize_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_index_resize_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_index_resize_1/index_resize_req
      -- CP-element group 35: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_index_resize_1/index_resize_ack
      -- CP-element group 35: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_index_scale_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_index_scale_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_index_scale_1/scale_rename_req
      -- CP-element group 35: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_index_scale_1/scale_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_final_index_sum_regn_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_final_index_sum_regn_Sample/req
      -- 
    ca_5776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2282_inst_ack_1, ack => convTransposeC_CP_5489_elements(35)); -- 
    req_5801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(35), ack => array_obj_ref_2288_index_offset_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	55 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_final_index_sum_regn_sample_complete
      -- CP-element group 36: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_final_index_sum_regn_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_final_index_sum_regn_Sample/ack
      -- 
    ack_5802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2288_index_offset_ack_0, ack => convTransposeC_CP_5489_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	89 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (11) 
      -- CP-element group 37: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2289_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_offset_calculated
      -- CP-element group 37: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_final_index_sum_regn_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_final_index_sum_regn_Update/ack
      -- CP-element group 37: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_base_plus_offset/$entry
      -- CP-element group 37: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_base_plus_offset/$exit
      -- CP-element group 37: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_base_plus_offset/sum_rename_req
      -- CP-element group 37: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2289_request/$entry
      -- CP-element group 37: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2289_request/req
      -- 
    ack_5807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2288_index_offset_ack_1, ack => convTransposeC_CP_5489_elements(37)); -- 
    req_5816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(37), ack => addr_of_2289_final_reg_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2289_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2289_request/$exit
      -- CP-element group 38: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2289_request/ack
      -- 
    ack_5817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2289_final_reg_ack_0, ack => convTransposeC_CP_5489_elements(38)); -- 
    -- CP-element group 39:  join  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	89 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (24) 
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2289_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2289_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2289_complete/ack
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_base_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_word_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_base_address_resized
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_base_addr_resize/$entry
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_base_addr_resize/$exit
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_base_addr_resize/base_resize_req
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_base_addr_resize/base_resize_ack
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_word_addrgen/$entry
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_word_addrgen/$exit
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_word_addrgen/root_register_req
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_word_addrgen/root_register_ack
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_Sample/word_access_start/$entry
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_Sample/word_access_start/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_Sample/word_access_start/word_0/rr
      -- 
    ack_5822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2289_final_reg_ack_1, ack => convTransposeC_CP_5489_elements(39)); -- 
    rr_5855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(39), ack => ptr_deref_2293_load_0_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_Sample/word_access_start/$exit
      -- CP-element group 40: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_Sample/word_access_start/word_0/$exit
      -- CP-element group 40: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_Sample/word_access_start/word_0/ra
      -- 
    ra_5856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2293_load_0_ack_0, ack => convTransposeC_CP_5489_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	89 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	50 
    -- CP-element group 41:  members (9) 
      -- CP-element group 41: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_Update/word_access_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_Update/word_access_complete/word_0/$exit
      -- CP-element group 41: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_Update/word_access_complete/word_0/ca
      -- CP-element group 41: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_Update/ptr_deref_2293_Merge/$entry
      -- CP-element group 41: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_Update/ptr_deref_2293_Merge/$exit
      -- CP-element group 41: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_Update/ptr_deref_2293_Merge/merge_req
      -- CP-element group 41: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_Update/ptr_deref_2293_Merge/merge_ack
      -- 
    ca_5867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2293_load_0_ack_1, ack => convTransposeC_CP_5489_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	89 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2298_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2298_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2298_Sample/ra
      -- 
    ra_5881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2298_inst_ack_0, ack => convTransposeC_CP_5489_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	89 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2298_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2298_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2298_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2312_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2312_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2312_Sample/rr
      -- 
    ca_5886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2298_inst_ack_1, ack => convTransposeC_CP_5489_elements(43)); -- 
    rr_5894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(43), ack => type_cast_2312_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2312_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2312_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2312_Sample/ra
      -- 
    ra_5895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2312_inst_ack_0, ack => convTransposeC_CP_5489_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	89 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (16) 
      -- CP-element group 45: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_index_scale_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_index_resize_1/index_resize_req
      -- CP-element group 45: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_index_scale_1/scale_rename_req
      -- CP-element group 45: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_index_scale_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_index_scale_1/scale_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_index_computed_1
      -- CP-element group 45: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_index_resize_1/index_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_index_resize_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_index_resize_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_final_index_sum_regn_Sample/req
      -- CP-element group 45: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_final_index_sum_regn_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2312_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2312_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2312_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_index_resized_1
      -- CP-element group 45: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_index_scaled_1
      -- 
    ca_5900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2312_inst_ack_1, ack => convTransposeC_CP_5489_elements(45)); -- 
    req_5925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(45), ack => array_obj_ref_2318_index_offset_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	55 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_final_index_sum_regn_sample_complete
      -- CP-element group 46: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_final_index_sum_regn_Sample/ack
      -- CP-element group 46: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_final_index_sum_regn_Sample/$exit
      -- 
    ack_5926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2318_index_offset_ack_0, ack => convTransposeC_CP_5489_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	89 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (11) 
      -- CP-element group 47: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_base_plus_offset/$entry
      -- CP-element group 47: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_final_index_sum_regn_Update/ack
      -- CP-element group 47: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_final_index_sum_regn_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2319_request/req
      -- CP-element group 47: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2319_request/$entry
      -- CP-element group 47: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_base_plus_offset/sum_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_base_plus_offset/sum_rename_req
      -- CP-element group 47: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_base_plus_offset/$exit
      -- CP-element group 47: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2319_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_root_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_offset_calculated
      -- 
    ack_5931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2318_index_offset_ack_1, ack => convTransposeC_CP_5489_elements(47)); -- 
    req_5940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(47), ack => addr_of_2319_final_reg_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2319_request/ack
      -- CP-element group 48: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2319_request/$exit
      -- CP-element group 48: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2319_sample_completed_
      -- 
    ack_5941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2319_final_reg_ack_0, ack => convTransposeC_CP_5489_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	89 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (19) 
      -- CP-element group 49: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_word_addrgen/root_register_req
      -- CP-element group 49: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_word_addrgen/root_register_ack
      -- CP-element group 49: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_base_addr_resize/base_resize_req
      -- CP-element group 49: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_base_addr_resize/base_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_base_addr_resize/$entry
      -- CP-element group 49: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_word_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_word_addrgen/$exit
      -- CP-element group 49: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_base_addr_resize/$exit
      -- CP-element group 49: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_word_addrgen/$entry
      -- CP-element group 49: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_base_address_resized
      -- CP-element group 49: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_base_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2319_complete/ack
      -- CP-element group 49: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2319_complete/$exit
      -- CP-element group 49: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2319_update_completed_
      -- 
    ack_5946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2319_final_reg_ack_1, ack => convTransposeC_CP_5489_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	41 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_Sample/ptr_deref_2322_Split/$entry
      -- CP-element group 50: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_Sample/ptr_deref_2322_Split/$exit
      -- CP-element group 50: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_Sample/ptr_deref_2322_Split/split_req
      -- CP-element group 50: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_Sample/word_access_start/word_0/rr
      -- CP-element group 50: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_Sample/word_access_start/word_0/$entry
      -- CP-element group 50: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_Sample/word_access_start/$entry
      -- CP-element group 50: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_Sample/ptr_deref_2322_Split/split_ack
      -- 
    rr_5984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(50), ack => ptr_deref_2322_store_0_req_0); -- 
    convTransposeC_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5489_elements(41) & convTransposeC_CP_5489_elements(49);
      gj_convTransposeC_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5489_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_Sample/word_access_start/word_0/ra
      -- CP-element group 51: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_Sample/word_access_start/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_Sample/word_access_start/$exit
      -- 
    ra_5985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2322_store_0_ack_0, ack => convTransposeC_CP_5489_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	89 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_Update/word_access_complete/word_0/ca
      -- CP-element group 52: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_Update/word_access_complete/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_Update/word_access_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_Update/$exit
      -- 
    ca_5996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2322_store_0_ack_1, ack => convTransposeC_CP_5489_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	89 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2328_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2328_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2328_sample_completed_
      -- 
    ra_6005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2328_inst_ack_0, ack => convTransposeC_CP_5489_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	89 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2328_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2328_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2328_update_completed_
      -- 
    ca_6010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2328_inst_ack_1, ack => convTransposeC_CP_5489_elements(54)); -- 
    -- CP-element group 55:  branch  join  transition  place  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	36 
    -- CP-element group 55: 	46 
    -- CP-element group 55: 	52 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (10) 
      -- CP-element group 55: 	 branch_block_stmt_2089/if_stmt_2343_dead_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_2089/if_stmt_2343_eval_test/$exit
      -- CP-element group 55: 	 branch_block_stmt_2089/if_stmt_2343_eval_test/branch_req
      -- CP-element group 55: 	 branch_block_stmt_2089/if_stmt_2343_if_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_2089/if_stmt_2343_eval_test/$entry
      -- CP-element group 55: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342__exit__
      -- CP-element group 55: 	 branch_block_stmt_2089/if_stmt_2343__entry__
      -- CP-element group 55: 	 branch_block_stmt_2089/R_cmp_2344_place
      -- CP-element group 55: 	 branch_block_stmt_2089/if_stmt_2343_else_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/$exit
      -- 
    branch_req_6018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(55), ack => if_stmt_2343_branch_req_0); -- 
    convTransposeC_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5489_elements(36) & convTransposeC_CP_5489_elements(46) & convTransposeC_CP_5489_elements(52) & convTransposeC_CP_5489_elements(54);
      gj_convTransposeC_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5489_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	84 
    -- CP-element group 56: 	85 
    -- CP-element group 56:  members (24) 
      -- CP-element group 56: 	 branch_block_stmt_2089/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2241/phi_stmt_2241_sources/type_cast_2244/SplitProtocol/Update/cr
      -- CP-element group 56: 	 branch_block_stmt_2089/merge_stmt_2349_PhiReqMerge
      -- CP-element group 56: 	 branch_block_stmt_2089/assign_stmt_2355/$entry
      -- CP-element group 56: 	 branch_block_stmt_2089/assign_stmt_2355/$exit
      -- CP-element group 56: 	 branch_block_stmt_2089/if_stmt_2343_if_link/if_choice_transition
      -- CP-element group 56: 	 branch_block_stmt_2089/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2241/phi_stmt_2241_sources/type_cast_2244/SplitProtocol/Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_2089/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_2089/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_2089/if_stmt_2343_if_link/$exit
      -- CP-element group 56: 	 branch_block_stmt_2089/assign_stmt_2355__entry__
      -- CP-element group 56: 	 branch_block_stmt_2089/merge_stmt_2349__exit__
      -- CP-element group 56: 	 branch_block_stmt_2089/ifx_xthen_whilex_xbody
      -- CP-element group 56: 	 branch_block_stmt_2089/assign_stmt_2355__exit__
      -- CP-element group 56: 	 branch_block_stmt_2089/whilex_xbody_ifx_xthen
      -- CP-element group 56: 	 branch_block_stmt_2089/merge_stmt_2349_PhiAck/$entry
      -- CP-element group 56: 	 branch_block_stmt_2089/merge_stmt_2349_PhiAck/$exit
      -- CP-element group 56: 	 branch_block_stmt_2089/merge_stmt_2349_PhiAck/dummy
      -- CP-element group 56: 	 branch_block_stmt_2089/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2241/phi_stmt_2241_sources/type_cast_2244/SplitProtocol/Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_2089/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2241/phi_stmt_2241_sources/type_cast_2244/SplitProtocol/Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_2089/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2241/phi_stmt_2241_sources/type_cast_2244/SplitProtocol/$entry
      -- CP-element group 56: 	 branch_block_stmt_2089/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2241/phi_stmt_2241_sources/type_cast_2244/$entry
      -- CP-element group 56: 	 branch_block_stmt_2089/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2241/phi_stmt_2241_sources/$entry
      -- CP-element group 56: 	 branch_block_stmt_2089/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2241/$entry
      -- CP-element group 56: 	 branch_block_stmt_2089/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- 
    if_choice_transition_6023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2343_branch_ack_1, ack => convTransposeC_CP_5489_elements(56)); -- 
    cr_6226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(56), ack => type_cast_2244_inst_req_1); -- 
    rr_6221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(56), ack => type_cast_2244_inst_req_0); -- 
    -- CP-element group 57:  fork  transition  place  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	59 
    -- CP-element group 57: 	61 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (24) 
      -- CP-element group 57: 	 branch_block_stmt_2089/merge_stmt_2357_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_2089/merge_stmt_2357_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_2089/merge_stmt_2357_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_2089/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/$entry
      -- CP-element group 57: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2393_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2367_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_2089/if_stmt_2343_else_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_2089/merge_stmt_2357_PhiAck/dummy
      -- CP-element group 57: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2393_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2393_update_start_
      -- CP-element group 57: 	 branch_block_stmt_2089/if_stmt_2343_else_link/else_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_2089/merge_stmt_2357__exit__
      -- CP-element group 57: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399__entry__
      -- CP-element group 57: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2376_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_2089/whilex_xbody_ifx_xelse
      -- CP-element group 57: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2376_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2376_update_start_
      -- CP-element group 57: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2367_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2367_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2367_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2367_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2367_update_start_
      -- CP-element group 57: 	 branch_block_stmt_2089/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- 
    else_choice_transition_6027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2343_branch_ack_0, ack => convTransposeC_CP_5489_elements(57)); -- 
    cr_6076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(57), ack => type_cast_2393_inst_req_1); -- 
    cr_6062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(57), ack => type_cast_2376_inst_req_1); -- 
    cr_6048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(57), ack => type_cast_2367_inst_req_1); -- 
    rr_6043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(57), ack => type_cast_2367_inst_req_0); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2367_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2367_Sample/ra
      -- CP-element group 58: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2367_Sample/$exit
      -- 
    ra_6044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2367_inst_ack_0, ack => convTransposeC_CP_5489_elements(58)); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2376_Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2376_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2376_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2367_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2367_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2367_update_completed_
      -- 
    ca_6049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2367_inst_ack_1, ack => convTransposeC_CP_5489_elements(59)); -- 
    rr_6057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(59), ack => type_cast_2376_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2376_Sample/ra
      -- CP-element group 60: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2376_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2376_sample_completed_
      -- 
    ra_6058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2376_inst_ack_0, ack => convTransposeC_CP_5489_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	57 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2393_Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2376_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2393_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2376_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2393_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2376_update_completed_
      -- 
    ca_6063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2376_inst_ack_1, ack => convTransposeC_CP_5489_elements(61)); -- 
    rr_6071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(61), ack => type_cast_2393_inst_req_0); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2393_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2393_Sample/ra
      -- CP-element group 62: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2393_sample_completed_
      -- 
    ra_6072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2393_inst_ack_0, ack => convTransposeC_CP_5489_elements(62)); -- 
    -- CP-element group 63:  branch  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (13) 
      -- CP-element group 63: 	 branch_block_stmt_2089/if_stmt_2400_if_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_2089/if_stmt_2400_eval_test/branch_req
      -- CP-element group 63: 	 branch_block_stmt_2089/if_stmt_2400_eval_test/$entry
      -- CP-element group 63: 	 branch_block_stmt_2089/if_stmt_2400_eval_test/$exit
      -- CP-element group 63: 	 branch_block_stmt_2089/R_cmp128_2401_place
      -- CP-element group 63: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2393_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_2089/if_stmt_2400_else_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/$exit
      -- CP-element group 63: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2393_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399/type_cast_2393_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_2089/if_stmt_2400_dead_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_2089/assign_stmt_2363_to_assign_stmt_2399__exit__
      -- CP-element group 63: 	 branch_block_stmt_2089/if_stmt_2400__entry__
      -- 
    ca_6077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2393_inst_ack_1, ack => convTransposeC_CP_5489_elements(63)); -- 
    branch_req_6085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(63), ack => if_stmt_2400_branch_req_0); -- 
    -- CP-element group 64:  merge  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (15) 
      -- CP-element group 64: 	 branch_block_stmt_2089/if_stmt_2400_if_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_2089/if_stmt_2400_if_link/if_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_2089/merge_stmt_2406_PhiReqMerge
      -- CP-element group 64: 	 branch_block_stmt_2089/ifx_xelse_whilex_xend
      -- CP-element group 64: 	 branch_block_stmt_2089/assign_stmt_2411/$entry
      -- CP-element group 64: 	 branch_block_stmt_2089/assign_stmt_2411/WPIPE_Block2_done_2408_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_2089/assign_stmt_2411/WPIPE_Block2_done_2408_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_2089/assign_stmt_2411/WPIPE_Block2_done_2408_Sample/req
      -- CP-element group 64: 	 branch_block_stmt_2089/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_2089/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 64: 	 branch_block_stmt_2089/merge_stmt_2406__exit__
      -- CP-element group 64: 	 branch_block_stmt_2089/assign_stmt_2411__entry__
      -- CP-element group 64: 	 branch_block_stmt_2089/merge_stmt_2406_PhiAck/$entry
      -- CP-element group 64: 	 branch_block_stmt_2089/merge_stmt_2406_PhiAck/$exit
      -- CP-element group 64: 	 branch_block_stmt_2089/merge_stmt_2406_PhiAck/dummy
      -- 
    if_choice_transition_6090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2400_branch_ack_1, ack => convTransposeC_CP_5489_elements(64)); -- 
    req_6107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(64), ack => WPIPE_Block2_done_2408_inst_req_0); -- 
    -- CP-element group 65:  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	73 
    -- CP-element group 65: 	74 
    -- CP-element group 65: 	76 
    -- CP-element group 65: 	77 
    -- CP-element group 65:  members (20) 
      -- CP-element group 65: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/$entry
      -- CP-element group 65: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/$entry
      -- CP-element group 65: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 65: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_2089/if_stmt_2400_else_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_2089/if_stmt_2400_else_link/else_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/SplitProtocol/Update/cr
      -- CP-element group 65: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/$entry
      -- CP-element group 65: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/SplitProtocol/Update/cr
      -- CP-element group 65: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/$entry
      -- CP-element group 65: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/$entry
      -- 
    else_choice_transition_6094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2400_branch_ack_0, ack => convTransposeC_CP_5489_elements(65)); -- 
    rr_6166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(65), ack => type_cast_2187_inst_req_0); -- 
    cr_6171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(65), ack => type_cast_2187_inst_req_1); -- 
    cr_6194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(65), ack => type_cast_2181_inst_req_1); -- 
    rr_6189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(65), ack => type_cast_2181_inst_req_0); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_2089/assign_stmt_2411/WPIPE_Block2_done_2408_Update/req
      -- CP-element group 66: 	 branch_block_stmt_2089/assign_stmt_2411/WPIPE_Block2_done_2408_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_2089/assign_stmt_2411/WPIPE_Block2_done_2408_update_start_
      -- CP-element group 66: 	 branch_block_stmt_2089/assign_stmt_2411/WPIPE_Block2_done_2408_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_2089/assign_stmt_2411/WPIPE_Block2_done_2408_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_2089/assign_stmt_2411/WPIPE_Block2_done_2408_Sample/ack
      -- 
    ack_6108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2408_inst_ack_0, ack => convTransposeC_CP_5489_elements(66)); -- 
    req_6112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(66), ack => WPIPE_Block2_done_2408_inst_req_1); -- 
    -- CP-element group 67:  transition  place  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (16) 
      -- CP-element group 67: 	 branch_block_stmt_2089/assign_stmt_2411/WPIPE_Block2_done_2408_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_2089/merge_stmt_2413_PhiReqMerge
      -- CP-element group 67: 	 $exit
      -- CP-element group 67: 	 branch_block_stmt_2089/assign_stmt_2411/$exit
      -- CP-element group 67: 	 branch_block_stmt_2089/branch_block_stmt_2089__exit__
      -- CP-element group 67: 	 branch_block_stmt_2089/assign_stmt_2411/WPIPE_Block2_done_2408_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_2089/assign_stmt_2411/WPIPE_Block2_done_2408_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_2089/$exit
      -- CP-element group 67: 	 branch_block_stmt_2089/merge_stmt_2413__exit__
      -- CP-element group 67: 	 branch_block_stmt_2089/assign_stmt_2411__exit__
      -- CP-element group 67: 	 branch_block_stmt_2089/return__
      -- CP-element group 67: 	 branch_block_stmt_2089/return___PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2089/return___PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_2089/merge_stmt_2413_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_2089/merge_stmt_2413_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_2089/merge_stmt_2413_PhiAck/dummy
      -- 
    ack_6113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2408_inst_ack_1, ack => convTransposeC_CP_5489_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	31 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/SplitProtocol/Sample/ra
      -- CP-element group 68: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/SplitProtocol/Sample/$exit
      -- 
    ra_6133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2185_inst_ack_0, ack => convTransposeC_CP_5489_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	31 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/SplitProtocol/Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/SplitProtocol/Update/ca
      -- 
    ca_6138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2185_inst_ack_1, ack => convTransposeC_CP_5489_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (5) 
      -- CP-element group 70: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/$exit
      -- CP-element group 70: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_req
      -- CP-element group 70: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/$exit
      -- CP-element group 70: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/$exit
      -- CP-element group 70: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2185/SplitProtocol/$exit
      -- 
    phi_stmt_2182_req_6139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2182_req_6139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(70), ack => phi_stmt_2182_req_0); -- 
    convTransposeC_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5489_elements(68) & convTransposeC_CP_5489_elements(69);
      gj_convTransposeC_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5489_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  transition  output  delay-element  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	31 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/$exit
      -- CP-element group 71: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/phi_stmt_2175_req
      -- CP-element group 71: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2179_konst_delay_trans
      -- CP-element group 71: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/$exit
      -- 
    phi_stmt_2175_req_6147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2175_req_6147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(71), ack => phi_stmt_2175_req_0); -- 
    -- Element group convTransposeC_CP_5489_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => convTransposeC_CP_5489_elements(31), ack => convTransposeC_CP_5489_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  join  transition  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	80 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_2089/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5489_elements(70) & convTransposeC_CP_5489_elements(71);
      gj_convTransposeC_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5489_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	65 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/SplitProtocol/Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/SplitProtocol/Sample/ra
      -- 
    ra_6167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2187_inst_ack_0, ack => convTransposeC_CP_5489_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	65 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/SplitProtocol/Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/SplitProtocol/Update/ca
      -- 
    ca_6172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2187_inst_ack_1, ack => convTransposeC_CP_5489_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	79 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/$exit
      -- CP-element group 75: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_req
      -- CP-element group 75: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/$exit
      -- CP-element group 75: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/SplitProtocol/$exit
      -- CP-element group 75: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2182/phi_stmt_2182_sources/type_cast_2187/$exit
      -- 
    phi_stmt_2182_req_6173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2182_req_6173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(75), ack => phi_stmt_2182_req_1); -- 
    convTransposeC_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5489_elements(73) & convTransposeC_CP_5489_elements(74);
      gj_convTransposeC_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5489_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	65 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/SplitProtocol/Sample/ra
      -- CP-element group 76: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/SplitProtocol/Sample/$exit
      -- 
    ra_6190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2181_inst_ack_0, ack => convTransposeC_CP_5489_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	65 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/SplitProtocol/Update/ca
      -- CP-element group 77: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/SplitProtocol/Update/$exit
      -- 
    ca_6195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2181_inst_ack_1, ack => convTransposeC_CP_5489_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/$exit
      -- CP-element group 78: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/phi_stmt_2175_req
      -- CP-element group 78: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/SplitProtocol/$exit
      -- CP-element group 78: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/$exit
      -- CP-element group 78: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/$exit
      -- 
    phi_stmt_2175_req_6196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2175_req_6196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(78), ack => phi_stmt_2175_req_1); -- 
    convTransposeC_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5489_elements(76) & convTransposeC_CP_5489_elements(77);
      gj_convTransposeC_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5489_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	75 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_2089/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5489_elements(75) & convTransposeC_CP_5489_elements(78);
      gj_convTransposeC_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5489_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  merge  fork  transition  place  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	72 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_2089/merge_stmt_2174_PhiReqMerge
      -- CP-element group 80: 	 branch_block_stmt_2089/merge_stmt_2174_PhiAck/$entry
      -- 
    convTransposeC_CP_5489_elements(80) <= OrReduce(convTransposeC_CP_5489_elements(72) & convTransposeC_CP_5489_elements(79));
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2089/merge_stmt_2174_PhiAck/phi_stmt_2175_ack
      -- 
    phi_stmt_2175_ack_6201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2175_ack_0, ack => convTransposeC_CP_5489_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_2089/merge_stmt_2174_PhiAck/phi_stmt_2182_ack
      -- 
    phi_stmt_2182_ack_6202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2182_ack_0, ack => convTransposeC_CP_5489_elements(82)); -- 
    -- CP-element group 83:  join  transition  place  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	87 
    -- CP-element group 83:  members (10) 
      -- CP-element group 83: 	 branch_block_stmt_2089/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 83: 	 branch_block_stmt_2089/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2241/$entry
      -- CP-element group 83: 	 branch_block_stmt_2089/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2241/phi_stmt_2241_sources/$entry
      -- CP-element group 83: 	 branch_block_stmt_2089/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 83: 	 branch_block_stmt_2089/assign_stmt_2193_to_assign_stmt_2238__exit__
      -- CP-element group 83: 	 branch_block_stmt_2089/merge_stmt_2174__exit__
      -- CP-element group 83: 	 branch_block_stmt_2089/assign_stmt_2193_to_assign_stmt_2238__entry__
      -- CP-element group 83: 	 branch_block_stmt_2089/merge_stmt_2174_PhiAck/$exit
      -- CP-element group 83: 	 branch_block_stmt_2089/assign_stmt_2193_to_assign_stmt_2238/$entry
      -- CP-element group 83: 	 branch_block_stmt_2089/assign_stmt_2193_to_assign_stmt_2238/$exit
      -- 
    convTransposeC_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5489_elements(81) & convTransposeC_CP_5489_elements(82);
      gj_convTransposeC_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5489_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	56 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_2089/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2241/phi_stmt_2241_sources/type_cast_2244/SplitProtocol/Sample/ra
      -- CP-element group 84: 	 branch_block_stmt_2089/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2241/phi_stmt_2241_sources/type_cast_2244/SplitProtocol/Sample/$exit
      -- 
    ra_6222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2244_inst_ack_0, ack => convTransposeC_CP_5489_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	56 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_2089/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2241/phi_stmt_2241_sources/type_cast_2244/SplitProtocol/Update/ca
      -- CP-element group 85: 	 branch_block_stmt_2089/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2241/phi_stmt_2241_sources/type_cast_2244/SplitProtocol/Update/$exit
      -- 
    ca_6227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2244_inst_ack_1, ack => convTransposeC_CP_5489_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_2089/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2241/phi_stmt_2241_req
      -- CP-element group 86: 	 branch_block_stmt_2089/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2241/phi_stmt_2241_sources/type_cast_2244/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_2089/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2241/phi_stmt_2241_sources/type_cast_2244/$exit
      -- CP-element group 86: 	 branch_block_stmt_2089/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2241/phi_stmt_2241_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_2089/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2241/$exit
      -- CP-element group 86: 	 branch_block_stmt_2089/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- 
    phi_stmt_2241_req_6228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2241_req_6228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(86), ack => phi_stmt_2241_req_0); -- 
    convTransposeC_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5489_elements(84) & convTransposeC_CP_5489_elements(85);
      gj_convTransposeC_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5489_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  output  delay-element  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	83 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_2089/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 87: 	 branch_block_stmt_2089/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2241/$exit
      -- CP-element group 87: 	 branch_block_stmt_2089/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2241/phi_stmt_2241_sources/$exit
      -- CP-element group 87: 	 branch_block_stmt_2089/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2241/phi_stmt_2241_sources/type_cast_2247_konst_delay_trans
      -- CP-element group 87: 	 branch_block_stmt_2089/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2241/phi_stmt_2241_req
      -- 
    phi_stmt_2241_req_6239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2241_req_6239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(87), ack => phi_stmt_2241_req_1); -- 
    -- Element group convTransposeC_CP_5489_elements(87) is a control-delay.
    cp_element_87_delay: control_delay_element  generic map(name => " 87_delay", delay_value => 1)  port map(req => convTransposeC_CP_5489_elements(83), ack => convTransposeC_CP_5489_elements(87), clk => clk, reset =>reset);
    -- CP-element group 88:  merge  transition  place  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_2089/merge_stmt_2240_PhiReqMerge
      -- CP-element group 88: 	 branch_block_stmt_2089/merge_stmt_2240_PhiAck/$entry
      -- 
    convTransposeC_CP_5489_elements(88) <= OrReduce(convTransposeC_CP_5489_elements(86) & convTransposeC_CP_5489_elements(87));
    -- CP-element group 89:  fork  transition  place  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	37 
    -- CP-element group 89: 	39 
    -- CP-element group 89: 	41 
    -- CP-element group 89: 	42 
    -- CP-element group 89: 	43 
    -- CP-element group 89: 	45 
    -- CP-element group 89: 	47 
    -- CP-element group 89: 	49 
    -- CP-element group 89: 	52 
    -- CP-element group 89: 	53 
    -- CP-element group 89: 	54 
    -- CP-element group 89: 	32 
    -- CP-element group 89: 	33 
    -- CP-element group 89: 	35 
    -- CP-element group 89:  members (51) 
      -- CP-element group 89: 	 branch_block_stmt_2089/merge_stmt_2240_PhiAck/$exit
      -- CP-element group 89: 	 branch_block_stmt_2089/merge_stmt_2240_PhiAck/phi_stmt_2241_ack
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2328_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_final_index_sum_regn_Update/req
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_final_index_sum_regn_update_start
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2318_final_index_sum_regn_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_2089/merge_stmt_2240__exit__
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342__entry__
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2328_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2328_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_update_start_
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2328_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2328_update_start_
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2328_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_Update/word_access_complete/word_0/cr
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2319_complete/req
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_Update/word_access_complete/word_0/$entry
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2319_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_Update/word_access_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2322_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/$entry
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2268_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2268_update_start_
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2268_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2268_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2268_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2268_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2282_update_start_
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2282_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2282_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2289_update_start_
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_final_index_sum_regn_update_start
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_final_index_sum_regn_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/array_obj_ref_2288_final_index_sum_regn_Update/req
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2289_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2289_complete/req
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_update_start_
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_Update/word_access_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_Update/word_access_complete/word_0/$entry
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/ptr_deref_2293_Update/word_access_complete/word_0/cr
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2298_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2298_update_start_
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2298_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2298_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2298_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2298_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2312_update_start_
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2312_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/type_cast_2312_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_2089/assign_stmt_2254_to_assign_stmt_2342/addr_of_2319_update_start_
      -- 
    phi_stmt_2241_ack_6244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2241_ack_0, ack => convTransposeC_CP_5489_elements(89)); -- 
    cr_6009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(89), ack => type_cast_2328_inst_req_1); -- 
    req_5930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(89), ack => array_obj_ref_2318_index_offset_req_1); -- 
    rr_6004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(89), ack => type_cast_2328_inst_req_0); -- 
    cr_5995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(89), ack => ptr_deref_2322_store_0_req_1); -- 
    req_5945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(89), ack => addr_of_2319_final_reg_req_1); -- 
    rr_5756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(89), ack => type_cast_2268_inst_req_0); -- 
    cr_5761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(89), ack => type_cast_2268_inst_req_1); -- 
    cr_5775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(89), ack => type_cast_2282_inst_req_1); -- 
    req_5806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(89), ack => array_obj_ref_2288_index_offset_req_1); -- 
    req_5821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(89), ack => addr_of_2289_final_reg_req_1); -- 
    cr_5866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(89), ack => ptr_deref_2293_load_0_req_1); -- 
    rr_5880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(89), ack => type_cast_2298_inst_req_0); -- 
    cr_5885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(89), ack => type_cast_2298_inst_req_1); -- 
    cr_5899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5489_elements(89), ack => type_cast_2312_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2276_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2306_wire : std_logic_vector(31 downto 0);
    signal R_idxprom97_2317_resized : std_logic_vector(13 downto 0);
    signal R_idxprom97_2317_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2287_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2287_scaled : std_logic_vector(13 downto 0);
    signal add102_2335 : std_logic_vector(31 downto 0);
    signal add44_2259 : std_logic_vector(15 downto 0);
    signal add88_2264 : std_logic_vector(15 downto 0);
    signal array_obj_ref_2288_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2288_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2288_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2288_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2288_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2288_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2318_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2318_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2318_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2318_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2318_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2318_root_address : std_logic_vector(13 downto 0);
    signal arrayidx92_2290 : std_logic_vector(31 downto 0);
    signal arrayidx98_2320 : std_logic_vector(31 downto 0);
    signal call11_2110 : std_logic_vector(15 downto 0);
    signal call13_2113 : std_logic_vector(15 downto 0);
    signal call14_2116 : std_logic_vector(15 downto 0);
    signal call15_2119 : std_logic_vector(15 downto 0);
    signal call17_2122 : std_logic_vector(15 downto 0);
    signal call19_2125 : std_logic_vector(15 downto 0);
    signal call1_2095 : std_logic_vector(15 downto 0);
    signal call3_2098 : std_logic_vector(15 downto 0);
    signal call5_2101 : std_logic_vector(15 downto 0);
    signal call7_2104 : std_logic_vector(15 downto 0);
    signal call9_2107 : std_logic_vector(15 downto 0);
    signal call_2092 : std_logic_vector(15 downto 0);
    signal cmp118_2373 : std_logic_vector(0 downto 0);
    signal cmp128_2399 : std_logic_vector(0 downto 0);
    signal cmp_2342 : std_logic_vector(0 downto 0);
    signal conv101_2329 : std_logic_vector(31 downto 0);
    signal conv105_2136 : std_logic_vector(31 downto 0);
    signal conv113_2368 : std_logic_vector(31 downto 0);
    signal conv116_2140 : std_logic_vector(31 downto 0);
    signal conv124_2394 : std_logic_vector(31 downto 0);
    signal conv127_2150 : std_logic_vector(31 downto 0);
    signal conv91_2269 : std_logic_vector(31 downto 0);
    signal conv95_2299 : std_logic_vector(31 downto 0);
    signal div117_2146 : std_logic_vector(31 downto 0);
    signal div_2132 : std_logic_vector(15 downto 0);
    signal idxprom97_2313 : std_logic_vector(63 downto 0);
    signal idxprom_2283 : std_logic_vector(63 downto 0);
    signal inc122_2377 : std_logic_vector(15 downto 0);
    signal inc122x_xinput_dim0x_x2_2382 : std_logic_vector(15 downto 0);
    signal inc_2363 : std_logic_vector(15 downto 0);
    signal indvar_2241 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2355 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2182 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2175 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2389 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2254 : std_logic_vector(15 downto 0);
    signal ptr_deref_2293_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2293_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2293_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2293_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2293_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2322_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2322_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2322_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2322_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2322_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2322_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr96_2308 : std_logic_vector(31 downto 0);
    signal shr_2278 : std_logic_vector(31 downto 0);
    signal tmp10_2238 : std_logic_vector(15 downto 0);
    signal tmp155_2193 : std_logic_vector(15 downto 0);
    signal tmp156_2198 : std_logic_vector(15 downto 0);
    signal tmp157_2203 : std_logic_vector(15 downto 0);
    signal tmp1_2161 : std_logic_vector(15 downto 0);
    signal tmp2_2208 : std_logic_vector(15 downto 0);
    signal tmp3_2213 : std_logic_vector(15 downto 0);
    signal tmp4_2167 : std_logic_vector(15 downto 0);
    signal tmp5_2172 : std_logic_vector(15 downto 0);
    signal tmp6_2218 : std_logic_vector(15 downto 0);
    signal tmp7_2223 : std_logic_vector(15 downto 0);
    signal tmp8_2228 : std_logic_vector(15 downto 0);
    signal tmp93_2294 : std_logic_vector(63 downto 0);
    signal tmp9_2233 : std_logic_vector(15 downto 0);
    signal tmp_2156 : std_logic_vector(15 downto 0);
    signal type_cast_2130_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2144_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2154_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2165_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2179_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2181_wire : std_logic_vector(15 downto 0);
    signal type_cast_2185_wire : std_logic_vector(15 downto 0);
    signal type_cast_2187_wire : std_logic_vector(15 downto 0);
    signal type_cast_2244_wire : std_logic_vector(15 downto 0);
    signal type_cast_2247_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2252_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2267_wire : std_logic_vector(31 downto 0);
    signal type_cast_2272_wire : std_logic_vector(31 downto 0);
    signal type_cast_2275_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2281_wire : std_logic_vector(63 downto 0);
    signal type_cast_2297_wire : std_logic_vector(31 downto 0);
    signal type_cast_2302_wire : std_logic_vector(31 downto 0);
    signal type_cast_2305_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2311_wire : std_logic_vector(63 downto 0);
    signal type_cast_2327_wire : std_logic_vector(31 downto 0);
    signal type_cast_2333_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2338_wire : std_logic_vector(31 downto 0);
    signal type_cast_2340_wire : std_logic_vector(31 downto 0);
    signal type_cast_2353_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2361_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2366_wire : std_logic_vector(31 downto 0);
    signal type_cast_2386_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2392_wire : std_logic_vector(31 downto 0);
    signal type_cast_2410_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2288_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2288_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2288_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2288_resized_base_address <= "00000000000000";
    array_obj_ref_2318_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2318_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2318_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2318_resized_base_address <= "00000000000000";
    ptr_deref_2293_word_offset_0 <= "00000000000000";
    ptr_deref_2322_word_offset_0 <= "00000000000000";
    type_cast_2130_wire_constant <= "0000000000000001";
    type_cast_2144_wire_constant <= "00000000000000000000000000000001";
    type_cast_2154_wire_constant <= "1111111111111111";
    type_cast_2165_wire_constant <= "1111111111111111";
    type_cast_2179_wire_constant <= "0000000000000000";
    type_cast_2247_wire_constant <= "0000000000000000";
    type_cast_2252_wire_constant <= "0000000000000100";
    type_cast_2275_wire_constant <= "00000000000000000000000000000010";
    type_cast_2305_wire_constant <= "00000000000000000000000000000010";
    type_cast_2333_wire_constant <= "00000000000000000000000000000100";
    type_cast_2353_wire_constant <= "0000000000000001";
    type_cast_2361_wire_constant <= "0000000000000001";
    type_cast_2386_wire_constant <= "0000000000000000";
    type_cast_2410_wire_constant <= "0000000000000001";
    phi_stmt_2175: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2179_wire_constant & type_cast_2181_wire;
      req <= phi_stmt_2175_req_0 & phi_stmt_2175_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2175",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2175_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2175,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2175
    phi_stmt_2182: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2185_wire & type_cast_2187_wire;
      req <= phi_stmt_2182_req_0 & phi_stmt_2182_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2182",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2182_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2182,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2182
    phi_stmt_2241: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2244_wire & type_cast_2247_wire_constant;
      req <= phi_stmt_2241_req_0 & phi_stmt_2241_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2241",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2241_ack_0,
          idata => idata,
          odata => indvar_2241,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2241
    -- flow-through select operator MUX_2388_inst
    input_dim1x_x2_2389 <= type_cast_2386_wire_constant when (cmp118_2373(0) /=  '0') else inc_2363;
    addr_of_2289_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2289_final_reg_req_0;
      addr_of_2289_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2289_final_reg_req_1;
      addr_of_2289_final_reg_ack_1<= rack(0);
      addr_of_2289_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2289_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2288_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx92_2290,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2319_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2319_final_reg_req_0;
      addr_of_2319_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2319_final_reg_req_1;
      addr_of_2319_final_reg_ack_1<= rack(0);
      addr_of_2319_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2319_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2318_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx98_2320,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2135_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2135_inst_req_0;
      type_cast_2135_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2135_inst_req_1;
      type_cast_2135_inst_ack_1<= rack(0);
      type_cast_2135_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2135_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2098,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv105_2136,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2139_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2139_inst_req_0;
      type_cast_2139_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2139_inst_req_1;
      type_cast_2139_inst_ack_1<= rack(0);
      type_cast_2139_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2139_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_2095,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_2140,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2149_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2149_inst_req_0;
      type_cast_2149_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2149_inst_req_1;
      type_cast_2149_inst_ack_1<= rack(0);
      type_cast_2149_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2149_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2092,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv127_2150,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2181_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2181_inst_req_0;
      type_cast_2181_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2181_inst_req_1;
      type_cast_2181_inst_ack_1<= rack(0);
      type_cast_2181_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2181_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2389,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2181_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2185_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2185_inst_req_0;
      type_cast_2185_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2185_inst_req_1;
      type_cast_2185_inst_ack_1<= rack(0);
      type_cast_2185_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2185_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2132,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2185_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2187_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2187_inst_req_0;
      type_cast_2187_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2187_inst_req_1;
      type_cast_2187_inst_ack_1<= rack(0);
      type_cast_2187_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2187_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc122x_xinput_dim0x_x2_2382,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2187_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2244_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2244_inst_req_0;
      type_cast_2244_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2244_inst_req_1;
      type_cast_2244_inst_ack_1<= rack(0);
      type_cast_2244_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2244_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2355,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2244_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2268_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2268_inst_req_0;
      type_cast_2268_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2268_inst_req_1;
      type_cast_2268_inst_ack_1<= rack(0);
      type_cast_2268_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2268_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2267_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv91_2269,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2272_inst
    process(conv91_2269) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv91_2269(31 downto 0);
      type_cast_2272_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2277_inst
    process(ASHR_i32_i32_2276_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2276_wire(31 downto 0);
      shr_2278 <= tmp_var; -- 
    end process;
    type_cast_2282_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2282_inst_req_0;
      type_cast_2282_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2282_inst_req_1;
      type_cast_2282_inst_ack_1<= rack(0);
      type_cast_2282_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2282_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2281_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2283,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2298_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2298_inst_req_0;
      type_cast_2298_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2298_inst_req_1;
      type_cast_2298_inst_ack_1<= rack(0);
      type_cast_2298_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2298_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2297_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_2299,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2302_inst
    process(conv95_2299) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv95_2299(31 downto 0);
      type_cast_2302_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2307_inst
    process(ASHR_i32_i32_2306_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2306_wire(31 downto 0);
      shr96_2308 <= tmp_var; -- 
    end process;
    type_cast_2312_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2312_inst_req_0;
      type_cast_2312_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2312_inst_req_1;
      type_cast_2312_inst_ack_1<= rack(0);
      type_cast_2312_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2312_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2311_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom97_2313,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2328_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2328_inst_req_0;
      type_cast_2328_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2328_inst_req_1;
      type_cast_2328_inst_ack_1<= rack(0);
      type_cast_2328_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2328_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2327_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv101_2329,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2338_inst
    process(add102_2335) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add102_2335(31 downto 0);
      type_cast_2338_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2340_inst
    process(conv105_2136) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv105_2136(31 downto 0);
      type_cast_2340_wire <= tmp_var; -- 
    end process;
    type_cast_2367_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2367_inst_req_0;
      type_cast_2367_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2367_inst_req_1;
      type_cast_2367_inst_ack_1<= rack(0);
      type_cast_2367_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2367_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2366_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_2368,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2376_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2376_inst_req_0;
      type_cast_2376_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2376_inst_req_1;
      type_cast_2376_inst_ack_1<= rack(0);
      type_cast_2376_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2376_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp118_2373,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc122_2377,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2393_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2393_inst_req_0;
      type_cast_2393_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2393_inst_req_1;
      type_cast_2393_inst_ack_1<= rack(0);
      type_cast_2393_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2393_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2392_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv124_2394,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2288_index_1_rename
    process(R_idxprom_2287_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2287_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2287_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2288_index_1_resize
    process(idxprom_2283) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2283;
      ov := iv(13 downto 0);
      R_idxprom_2287_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2288_root_address_inst
    process(array_obj_ref_2288_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2288_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2288_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2318_index_1_rename
    process(R_idxprom97_2317_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom97_2317_resized;
      ov(13 downto 0) := iv;
      R_idxprom97_2317_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2318_index_1_resize
    process(idxprom97_2313) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom97_2313;
      ov := iv(13 downto 0);
      R_idxprom97_2317_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2318_root_address_inst
    process(array_obj_ref_2318_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2318_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2318_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2293_addr_0
    process(ptr_deref_2293_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2293_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2293_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2293_base_resize
    process(arrayidx92_2290) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx92_2290;
      ov := iv(13 downto 0);
      ptr_deref_2293_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2293_gather_scatter
    process(ptr_deref_2293_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2293_data_0;
      ov(63 downto 0) := iv;
      tmp93_2294 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2293_root_address_inst
    process(ptr_deref_2293_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2293_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2293_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2322_addr_0
    process(ptr_deref_2322_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2322_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2322_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2322_base_resize
    process(arrayidx98_2320) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx98_2320;
      ov := iv(13 downto 0);
      ptr_deref_2322_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2322_gather_scatter
    process(tmp93_2294) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp93_2294;
      ov(63 downto 0) := iv;
      ptr_deref_2322_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2322_root_address_inst
    process(ptr_deref_2322_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2322_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2322_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2343_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2342;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2343_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2343_branch_req_0,
          ack0 => if_stmt_2343_branch_ack_0,
          ack1 => if_stmt_2343_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2400_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp128_2399;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2400_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2400_branch_req_0,
          ack0 => if_stmt_2400_branch_ack_0,
          ack1 => if_stmt_2400_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2155_inst
    process(call9_2107) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2107, type_cast_2154_wire_constant, tmp_var);
      tmp_2156 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2166_inst
    process(call7_2104) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2104, type_cast_2165_wire_constant, tmp_var);
      tmp4_2167 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2197_inst
    process(input_dim1x_x1x_xph_2175, tmp155_2193) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2175, tmp155_2193, tmp_var);
      tmp156_2198 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2212_inst
    process(tmp1_2161, tmp2_2208) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp1_2161, tmp2_2208, tmp_var);
      tmp3_2213 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2222_inst
    process(tmp5_2172, tmp6_2218) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp5_2172, tmp6_2218, tmp_var);
      tmp7_2223 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2232_inst
    process(tmp3_2213, tmp8_2228) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_2213, tmp8_2228, tmp_var);
      tmp9_2233 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2258_inst
    process(tmp157_2203, input_dim2x_x1_2254) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp157_2203, input_dim2x_x1_2254, tmp_var);
      add44_2259 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2263_inst
    process(tmp10_2238, input_dim2x_x1_2254) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp10_2238, input_dim2x_x1_2254, tmp_var);
      add88_2264 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2354_inst
    process(indvar_2241) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2241, type_cast_2353_wire_constant, tmp_var);
      indvarx_xnext_2355 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2362_inst
    process(input_dim1x_x1x_xph_2175) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2175, type_cast_2361_wire_constant, tmp_var);
      inc_2363 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2381_inst
    process(inc122_2377, input_dim0x_x2x_xph_2182) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc122_2377, input_dim0x_x2x_xph_2182, tmp_var);
      inc122x_xinput_dim0x_x2_2382 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2334_inst
    process(conv101_2329) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv101_2329, type_cast_2333_wire_constant, tmp_var);
      add102_2335 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2276_inst
    process(type_cast_2272_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2272_wire, type_cast_2275_wire_constant, tmp_var);
      ASHR_i32_i32_2276_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2306_inst
    process(type_cast_2302_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2302_wire, type_cast_2305_wire_constant, tmp_var);
      ASHR_i32_i32_2306_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2372_inst
    process(conv113_2368, div117_2146) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv113_2368, div117_2146, tmp_var);
      cmp118_2373 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2398_inst
    process(conv124_2394, conv127_2150) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv124_2394, conv127_2150, tmp_var);
      cmp128_2399 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2131_inst
    process(call_2092) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2092, type_cast_2130_wire_constant, tmp_var);
      div_2132 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2145_inst
    process(conv116_2140) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv116_2140, type_cast_2144_wire_constant, tmp_var);
      div117_2146 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2192_inst
    process(call1_2095, input_dim0x_x2x_xph_2182) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call1_2095, input_dim0x_x2x_xph_2182, tmp_var);
      tmp155_2193 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2202_inst
    process(call3_2098, tmp156_2198) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call3_2098, tmp156_2198, tmp_var);
      tmp157_2203 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2207_inst
    process(call13_2113, input_dim1x_x1x_xph_2175) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_2113, input_dim1x_x1x_xph_2175, tmp_var);
      tmp2_2208 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2217_inst
    process(call13_2113, input_dim0x_x2x_xph_2182) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_2113, input_dim0x_x2x_xph_2182, tmp_var);
      tmp6_2218 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2227_inst
    process(call17_2122, tmp7_2223) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call17_2122, tmp7_2223, tmp_var);
      tmp8_2228 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2237_inst
    process(call19_2125, tmp9_2233) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call19_2125, tmp9_2233, tmp_var);
      tmp10_2238 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2253_inst
    process(indvar_2241) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2241, type_cast_2252_wire_constant, tmp_var);
      input_dim2x_x1_2254 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2341_inst
    process(type_cast_2338_wire, type_cast_2340_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2338_wire, type_cast_2340_wire, tmp_var);
      cmp_2342 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2160_inst
    process(tmp_2156, call14_2116) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp_2156, call14_2116, tmp_var);
      tmp1_2161 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2171_inst
    process(tmp4_2167, call14_2116) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp4_2167, call14_2116, tmp_var);
      tmp5_2172 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_2288_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2287_scaled;
      array_obj_ref_2288_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2288_index_offset_req_0;
      array_obj_ref_2288_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2288_index_offset_req_1;
      array_obj_ref_2288_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_2318_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom97_2317_scaled;
      array_obj_ref_2318_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2318_index_offset_req_0;
      array_obj_ref_2318_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2318_index_offset_req_1;
      array_obj_ref_2318_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- unary operator type_cast_2267_inst
    process(add44_2259) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add44_2259, tmp_var);
      type_cast_2267_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2281_inst
    process(shr_2278) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2278, tmp_var);
      type_cast_2281_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2297_inst
    process(add88_2264) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add88_2264, tmp_var);
      type_cast_2297_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2311_inst
    process(shr96_2308) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr96_2308, tmp_var);
      type_cast_2311_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2327_inst
    process(input_dim2x_x1_2254) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_2254, tmp_var);
      type_cast_2327_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2366_inst
    process(inc_2363) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2363, tmp_var);
      type_cast_2366_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2392_inst
    process(inc122x_xinput_dim0x_x2_2382) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc122x_xinput_dim0x_x2_2382, tmp_var);
      type_cast_2392_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_2293_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2293_load_0_req_0;
      ptr_deref_2293_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2293_load_0_req_1;
      ptr_deref_2293_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2293_word_address_0;
      ptr_deref_2293_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2322_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2322_store_0_req_0;
      ptr_deref_2322_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2322_store_0_req_1;
      ptr_deref_2322_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2322_word_address_0;
      data_in <= ptr_deref_2322_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_start_2091_inst RPIPE_Block2_start_2094_inst RPIPE_Block2_start_2097_inst RPIPE_Block2_start_2100_inst RPIPE_Block2_start_2103_inst RPIPE_Block2_start_2106_inst RPIPE_Block2_start_2109_inst RPIPE_Block2_start_2112_inst RPIPE_Block2_start_2115_inst RPIPE_Block2_start_2118_inst RPIPE_Block2_start_2121_inst RPIPE_Block2_start_2124_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(191 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 11 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 11 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant outBUFs : IntegerArray(11 downto 0) := (11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      reqL_unguarded(11) <= RPIPE_Block2_start_2091_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block2_start_2094_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block2_start_2097_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block2_start_2100_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block2_start_2103_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block2_start_2106_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block2_start_2109_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block2_start_2112_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block2_start_2115_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block2_start_2118_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block2_start_2121_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block2_start_2124_inst_req_0;
      RPIPE_Block2_start_2091_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block2_start_2094_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block2_start_2097_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block2_start_2100_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block2_start_2103_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block2_start_2106_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block2_start_2109_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block2_start_2112_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block2_start_2115_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block2_start_2118_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block2_start_2121_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block2_start_2124_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(11) <= RPIPE_Block2_start_2091_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block2_start_2094_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block2_start_2097_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block2_start_2100_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block2_start_2103_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block2_start_2106_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block2_start_2109_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block2_start_2112_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block2_start_2115_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block2_start_2118_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block2_start_2121_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block2_start_2124_inst_req_1;
      RPIPE_Block2_start_2091_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block2_start_2094_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block2_start_2097_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block2_start_2100_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block2_start_2103_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block2_start_2106_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block2_start_2109_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block2_start_2112_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block2_start_2115_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block2_start_2118_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block2_start_2121_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block2_start_2124_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      call_2092 <= data_out(191 downto 176);
      call1_2095 <= data_out(175 downto 160);
      call3_2098 <= data_out(159 downto 144);
      call5_2101 <= data_out(143 downto 128);
      call7_2104 <= data_out(127 downto 112);
      call9_2107 <= data_out(111 downto 96);
      call11_2110 <= data_out(95 downto 80);
      call13_2113 <= data_out(79 downto 64);
      call14_2116 <= data_out(63 downto 48);
      call15_2119 <= data_out(47 downto 32);
      call17_2122 <= data_out(31 downto 16);
      call19_2125 <= data_out(15 downto 0);
      Block2_start_read_0_gI: SplitGuardInterface generic map(name => "Block2_start_read_0_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_start_read_0: InputPortRevised -- 
        generic map ( name => "Block2_start_read_0", data_width => 16,  num_reqs => 12,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_start_pipe_read_req(0),
          oack => Block2_start_pipe_read_ack(0),
          odata => Block2_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2408_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2408_inst_req_0;
      WPIPE_Block2_done_2408_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2408_inst_req_1;
      WPIPE_Block2_done_2408_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2410_wire_constant;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_6285_start: Boolean;
  signal convTransposeD_CP_6285_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block3_start_2449_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2449_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2440_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2449_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2443_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2446_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2437_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2446_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2437_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2446_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2443_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2449_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2440_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2440_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2437_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2446_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2443_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2437_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2440_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2443_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2419_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2419_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2419_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2419_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2422_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2422_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2422_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2422_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2425_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2425_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2425_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2425_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2428_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2428_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2428_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2428_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2431_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2431_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2431_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2431_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2434_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2434_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2434_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2434_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2452_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2452_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2452_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2452_inst_ack_1 : boolean;
  signal type_cast_2469_inst_req_0 : boolean;
  signal type_cast_2469_inst_ack_0 : boolean;
  signal type_cast_2469_inst_req_1 : boolean;
  signal type_cast_2469_inst_ack_1 : boolean;
  signal type_cast_2473_inst_req_0 : boolean;
  signal type_cast_2473_inst_ack_0 : boolean;
  signal type_cast_2473_inst_req_1 : boolean;
  signal type_cast_2473_inst_ack_1 : boolean;
  signal type_cast_2477_inst_req_0 : boolean;
  signal type_cast_2477_inst_ack_0 : boolean;
  signal type_cast_2477_inst_req_1 : boolean;
  signal type_cast_2477_inst_ack_1 : boolean;
  signal type_cast_2595_inst_req_0 : boolean;
  signal type_cast_2595_inst_ack_0 : boolean;
  signal type_cast_2595_inst_req_1 : boolean;
  signal type_cast_2595_inst_ack_1 : boolean;
  signal type_cast_2609_inst_req_0 : boolean;
  signal type_cast_2609_inst_ack_0 : boolean;
  signal type_cast_2609_inst_req_1 : boolean;
  signal type_cast_2609_inst_ack_1 : boolean;
  signal array_obj_ref_2615_index_offset_req_0 : boolean;
  signal array_obj_ref_2615_index_offset_ack_0 : boolean;
  signal array_obj_ref_2615_index_offset_req_1 : boolean;
  signal array_obj_ref_2615_index_offset_ack_1 : boolean;
  signal addr_of_2616_final_reg_req_0 : boolean;
  signal addr_of_2616_final_reg_ack_0 : boolean;
  signal addr_of_2616_final_reg_req_1 : boolean;
  signal addr_of_2616_final_reg_ack_1 : boolean;
  signal ptr_deref_2620_load_0_req_0 : boolean;
  signal ptr_deref_2620_load_0_ack_0 : boolean;
  signal ptr_deref_2620_load_0_req_1 : boolean;
  signal ptr_deref_2620_load_0_ack_1 : boolean;
  signal type_cast_2625_inst_req_0 : boolean;
  signal type_cast_2625_inst_ack_0 : boolean;
  signal type_cast_2625_inst_req_1 : boolean;
  signal type_cast_2625_inst_ack_1 : boolean;
  signal type_cast_2639_inst_req_0 : boolean;
  signal type_cast_2639_inst_ack_0 : boolean;
  signal type_cast_2639_inst_req_1 : boolean;
  signal type_cast_2639_inst_ack_1 : boolean;
  signal array_obj_ref_2645_index_offset_req_0 : boolean;
  signal array_obj_ref_2645_index_offset_ack_0 : boolean;
  signal array_obj_ref_2645_index_offset_req_1 : boolean;
  signal array_obj_ref_2645_index_offset_ack_1 : boolean;
  signal addr_of_2646_final_reg_req_0 : boolean;
  signal addr_of_2646_final_reg_ack_0 : boolean;
  signal addr_of_2646_final_reg_req_1 : boolean;
  signal addr_of_2646_final_reg_ack_1 : boolean;
  signal ptr_deref_2649_store_0_req_0 : boolean;
  signal ptr_deref_2649_store_0_ack_0 : boolean;
  signal ptr_deref_2649_store_0_req_1 : boolean;
  signal ptr_deref_2649_store_0_ack_1 : boolean;
  signal type_cast_2655_inst_req_0 : boolean;
  signal type_cast_2655_inst_ack_0 : boolean;
  signal type_cast_2655_inst_req_1 : boolean;
  signal type_cast_2655_inst_ack_1 : boolean;
  signal if_stmt_2670_branch_req_0 : boolean;
  signal if_stmt_2670_branch_ack_1 : boolean;
  signal if_stmt_2670_branch_ack_0 : boolean;
  signal type_cast_2694_inst_req_0 : boolean;
  signal type_cast_2694_inst_ack_0 : boolean;
  signal type_cast_2694_inst_req_1 : boolean;
  signal type_cast_2694_inst_ack_1 : boolean;
  signal type_cast_2709_inst_req_0 : boolean;
  signal type_cast_2709_inst_ack_0 : boolean;
  signal type_cast_2709_inst_req_1 : boolean;
  signal type_cast_2709_inst_ack_1 : boolean;
  signal type_cast_2719_inst_req_0 : boolean;
  signal type_cast_2719_inst_ack_0 : boolean;
  signal type_cast_2719_inst_req_1 : boolean;
  signal type_cast_2719_inst_ack_1 : boolean;
  signal if_stmt_2726_branch_req_0 : boolean;
  signal if_stmt_2726_branch_ack_1 : boolean;
  signal if_stmt_2726_branch_ack_0 : boolean;
  signal WPIPE_Block3_done_2734_inst_req_0 : boolean;
  signal WPIPE_Block3_done_2734_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_2734_inst_req_1 : boolean;
  signal WPIPE_Block3_done_2734_inst_ack_1 : boolean;
  signal type_cast_2508_inst_req_0 : boolean;
  signal type_cast_2508_inst_ack_0 : boolean;
  signal type_cast_2508_inst_req_1 : boolean;
  signal type_cast_2508_inst_ack_1 : boolean;
  signal phi_stmt_2503_req_1 : boolean;
  signal type_cast_2514_inst_req_0 : boolean;
  signal type_cast_2514_inst_ack_0 : boolean;
  signal type_cast_2514_inst_req_1 : boolean;
  signal type_cast_2514_inst_ack_1 : boolean;
  signal phi_stmt_2509_req_1 : boolean;
  signal type_cast_2506_inst_req_0 : boolean;
  signal type_cast_2506_inst_ack_0 : boolean;
  signal type_cast_2506_inst_req_1 : boolean;
  signal type_cast_2506_inst_ack_1 : boolean;
  signal phi_stmt_2503_req_0 : boolean;
  signal type_cast_2512_inst_req_0 : boolean;
  signal type_cast_2512_inst_ack_0 : boolean;
  signal type_cast_2512_inst_req_1 : boolean;
  signal type_cast_2512_inst_ack_1 : boolean;
  signal phi_stmt_2509_req_0 : boolean;
  signal phi_stmt_2503_ack_0 : boolean;
  signal phi_stmt_2509_ack_0 : boolean;
  signal type_cast_2571_inst_req_0 : boolean;
  signal type_cast_2571_inst_ack_0 : boolean;
  signal type_cast_2571_inst_req_1 : boolean;
  signal type_cast_2571_inst_ack_1 : boolean;
  signal phi_stmt_2568_req_0 : boolean;
  signal phi_stmt_2568_req_1 : boolean;
  signal phi_stmt_2568_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_6285_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6285_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_6285_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6285_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_6285: Block -- control-path 
    signal convTransposeD_CP_6285_elements: BooleanArray(91 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_6285_elements(0) <= convTransposeD_CP_6285_start;
    convTransposeD_CP_6285_symbol <= convTransposeD_CP_6285_elements(67);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2417/$entry
      -- CP-element group 0: 	 branch_block_stmt_2417/branch_block_stmt_2417__entry__
      -- CP-element group 0: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453__entry__
      -- CP-element group 0: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/$entry
      -- CP-element group 0: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2419_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2419_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2419_Sample/rr
      -- 
    rr_6333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(0), ack => RPIPE_Block3_start_2419_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2419_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2419_update_start_
      -- CP-element group 1: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2419_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2419_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2419_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2419_Update/cr
      -- 
    ra_6334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2419_inst_ack_0, ack => convTransposeD_CP_6285_elements(1)); -- 
    cr_6338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(1), ack => RPIPE_Block3_start_2419_inst_req_1); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2419_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2419_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2419_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2422_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2422_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2422_Sample/rr
      -- 
    ca_6339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2419_inst_ack_1, ack => convTransposeD_CP_6285_elements(2)); -- 
    rr_6347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(2), ack => RPIPE_Block3_start_2422_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2422_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2422_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2422_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2422_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2422_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2422_Update/cr
      -- 
    ra_6348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2422_inst_ack_0, ack => convTransposeD_CP_6285_elements(3)); -- 
    cr_6352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(3), ack => RPIPE_Block3_start_2422_inst_req_1); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2422_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2422_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2422_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2425_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2425_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2425_Sample/rr
      -- 
    ca_6353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2422_inst_ack_1, ack => convTransposeD_CP_6285_elements(4)); -- 
    rr_6361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(4), ack => RPIPE_Block3_start_2425_inst_req_0); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2425_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2425_update_start_
      -- CP-element group 5: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2425_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2425_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2425_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2425_Update/cr
      -- 
    ra_6362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2425_inst_ack_0, ack => convTransposeD_CP_6285_elements(5)); -- 
    cr_6366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(5), ack => RPIPE_Block3_start_2425_inst_req_1); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2425_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2425_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2425_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2428_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2428_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2428_Sample/rr
      -- 
    ca_6367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2425_inst_ack_1, ack => convTransposeD_CP_6285_elements(6)); -- 
    rr_6375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(6), ack => RPIPE_Block3_start_2428_inst_req_0); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2428_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2428_update_start_
      -- CP-element group 7: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2428_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2428_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2428_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2428_Update/cr
      -- 
    ra_6376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2428_inst_ack_0, ack => convTransposeD_CP_6285_elements(7)); -- 
    cr_6380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(7), ack => RPIPE_Block3_start_2428_inst_req_1); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2428_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2428_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2428_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2431_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2431_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2431_Sample/rr
      -- 
    ca_6381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2428_inst_ack_1, ack => convTransposeD_CP_6285_elements(8)); -- 
    rr_6389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(8), ack => RPIPE_Block3_start_2431_inst_req_0); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2431_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2431_update_start_
      -- CP-element group 9: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2431_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2431_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2431_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2431_Update/cr
      -- 
    ra_6390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2431_inst_ack_0, ack => convTransposeD_CP_6285_elements(9)); -- 
    cr_6394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(9), ack => RPIPE_Block3_start_2431_inst_req_1); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2431_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2431_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2431_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2434_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2434_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2434_Sample/rr
      -- 
    ca_6395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2431_inst_ack_1, ack => convTransposeD_CP_6285_elements(10)); -- 
    rr_6403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(10), ack => RPIPE_Block3_start_2434_inst_req_0); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2434_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2434_update_start_
      -- CP-element group 11: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2434_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2434_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2434_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2434_Update/cr
      -- 
    ra_6404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2434_inst_ack_0, ack => convTransposeD_CP_6285_elements(11)); -- 
    cr_6408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(11), ack => RPIPE_Block3_start_2434_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2437_Sample/rr
      -- CP-element group 12: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2434_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2434_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2434_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2437_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2437_Sample/$entry
      -- 
    ca_6409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2434_inst_ack_1, ack => convTransposeD_CP_6285_elements(12)); -- 
    rr_6417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(12), ack => RPIPE_Block3_start_2437_inst_req_0); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2437_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2437_Update/cr
      -- CP-element group 13: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2437_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2437_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2437_update_start_
      -- CP-element group 13: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2437_Sample/$exit
      -- 
    ra_6418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2437_inst_ack_0, ack => convTransposeD_CP_6285_elements(13)); -- 
    cr_6422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(13), ack => RPIPE_Block3_start_2437_inst_req_1); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2437_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2440_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2440_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2437_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2440_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2437_update_completed_
      -- 
    ca_6423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2437_inst_ack_1, ack => convTransposeD_CP_6285_elements(14)); -- 
    rr_6431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(14), ack => RPIPE_Block3_start_2440_inst_req_0); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2440_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2440_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2440_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2440_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2440_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2440_Update/$entry
      -- 
    ra_6432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2440_inst_ack_0, ack => convTransposeD_CP_6285_elements(15)); -- 
    cr_6436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(15), ack => RPIPE_Block3_start_2440_inst_req_1); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2443_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2440_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2443_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2443_Sample/rr
      -- CP-element group 16: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2440_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2440_Update/$exit
      -- 
    ca_6437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2440_inst_ack_1, ack => convTransposeD_CP_6285_elements(16)); -- 
    rr_6445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(16), ack => RPIPE_Block3_start_2443_inst_req_0); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2443_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2443_update_start_
      -- CP-element group 17: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2443_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2443_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2443_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2443_Update/cr
      -- 
    ra_6446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2443_inst_ack_0, ack => convTransposeD_CP_6285_elements(17)); -- 
    cr_6450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(17), ack => RPIPE_Block3_start_2443_inst_req_1); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2443_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2443_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2446_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2446_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2446_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2443_Update/$exit
      -- 
    ca_6451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2443_inst_ack_1, ack => convTransposeD_CP_6285_elements(18)); -- 
    rr_6459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(18), ack => RPIPE_Block3_start_2446_inst_req_0); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2446_Update/cr
      -- CP-element group 19: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2446_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2446_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2446_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2446_update_start_
      -- CP-element group 19: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2446_Update/$entry
      -- 
    ra_6460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2446_inst_ack_0, ack => convTransposeD_CP_6285_elements(19)); -- 
    cr_6464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(19), ack => RPIPE_Block3_start_2446_inst_req_1); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2449_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2446_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2449_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2449_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2446_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2446_Update/$exit
      -- 
    ca_6465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2446_inst_ack_1, ack => convTransposeD_CP_6285_elements(20)); -- 
    rr_6473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(20), ack => RPIPE_Block3_start_2449_inst_req_0); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2449_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2449_Update/cr
      -- CP-element group 21: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2449_update_start_
      -- CP-element group 21: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2449_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2449_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2449_Update/$entry
      -- 
    ra_6474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2449_inst_ack_0, ack => convTransposeD_CP_6285_elements(21)); -- 
    cr_6478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(21), ack => RPIPE_Block3_start_2449_inst_req_1); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2449_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2449_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2452_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2449_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2452_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2452_Sample/rr
      -- 
    ca_6479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2449_inst_ack_1, ack => convTransposeD_CP_6285_elements(22)); -- 
    rr_6487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(22), ack => RPIPE_Block3_start_2452_inst_req_0); -- 
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2452_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2452_update_start_
      -- CP-element group 23: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2452_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2452_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2452_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2452_Update/cr
      -- 
    ra_6488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2452_inst_ack_0, ack => convTransposeD_CP_6285_elements(23)); -- 
    cr_6492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(23), ack => RPIPE_Block3_start_2452_inst_req_1); -- 
    -- CP-element group 24:  fork  transition  place  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	27 
    -- CP-element group 24: 	28 
    -- CP-element group 24: 	29 
    -- CP-element group 24: 	30 
    -- CP-element group 24:  members (25) 
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453__exit__
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500__entry__
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/$exit
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2452_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2452_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2420_to_assign_stmt_2453/RPIPE_Block3_start_2452_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/$entry
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2469_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2469_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2469_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2469_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2469_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2469_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2473_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2473_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2473_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2473_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2473_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2473_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2477_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2477_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2477_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2477_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2477_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2477_Update/cr
      -- 
    ca_6493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2452_inst_ack_1, ack => convTransposeD_CP_6285_elements(24)); -- 
    rr_6504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(24), ack => type_cast_2469_inst_req_0); -- 
    cr_6509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(24), ack => type_cast_2469_inst_req_1); -- 
    rr_6518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(24), ack => type_cast_2473_inst_req_0); -- 
    cr_6523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(24), ack => type_cast_2473_inst_req_1); -- 
    rr_6532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(24), ack => type_cast_2477_inst_req_0); -- 
    cr_6537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(24), ack => type_cast_2477_inst_req_1); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2469_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2469_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2469_Sample/ra
      -- 
    ra_6505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2469_inst_ack_0, ack => convTransposeD_CP_6285_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2469_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2469_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2469_Update/ca
      -- 
    ca_6510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2469_inst_ack_1, ack => convTransposeD_CP_6285_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	24 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2473_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2473_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2473_Sample/ra
      -- 
    ra_6519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2473_inst_ack_0, ack => convTransposeD_CP_6285_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	24 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2473_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2473_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2473_Update/ca
      -- 
    ca_6524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2473_inst_ack_1, ack => convTransposeD_CP_6285_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	24 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2477_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2477_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2477_Sample/ra
      -- 
    ra_6533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2477_inst_ack_0, ack => convTransposeD_CP_6285_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	24 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2477_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2477_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/type_cast_2477_Update/ca
      -- 
    ca_6538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2477_inst_ack_1, ack => convTransposeD_CP_6285_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	68 
    -- CP-element group 31: 	69 
    -- CP-element group 31: 	71 
    -- CP-element group 31: 	72 
    -- CP-element group 31:  members (20) 
      -- CP-element group 31: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500__exit__
      -- CP-element group 31: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_2417/assign_stmt_2460_to_assign_stmt_2500/$exit
      -- CP-element group 31: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/$entry
      -- CP-element group 31: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/$entry
      -- CP-element group 31: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Update/cr
      -- CP-element group 31: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/$entry
      -- CP-element group 31: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2514/$entry
      -- CP-element group 31: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2514/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2514/SplitProtocol/Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2514/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2514/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2514/SplitProtocol/Update/cr
      -- 
    rr_6928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(31), ack => type_cast_2508_inst_req_0); -- 
    cr_6933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(31), ack => type_cast_2508_inst_req_1); -- 
    rr_6951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(31), ack => type_cast_2514_inst_req_0); -- 
    cr_6956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(31), ack => type_cast_2514_inst_req_1); -- 
    convTransposeD_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6285_elements(26) & convTransposeD_CP_6285_elements(28) & convTransposeD_CP_6285_elements(30);
      gj_convTransposeD_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6285_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	91 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2595_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2595_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2595_Sample/ra
      -- 
    ra_6553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2595_inst_ack_0, ack => convTransposeD_CP_6285_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	91 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2595_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2595_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2595_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2609_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2609_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2609_Sample/rr
      -- 
    ca_6558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2595_inst_ack_1, ack => convTransposeD_CP_6285_elements(33)); -- 
    rr_6566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(33), ack => type_cast_2609_inst_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2609_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2609_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2609_Sample/ra
      -- 
    ra_6567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2609_inst_ack_0, ack => convTransposeD_CP_6285_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	91 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (16) 
      -- CP-element group 35: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2609_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2609_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2609_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_index_resized_1
      -- CP-element group 35: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_index_scaled_1
      -- CP-element group 35: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_index_computed_1
      -- CP-element group 35: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_index_resize_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_index_resize_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_index_resize_1/index_resize_req
      -- CP-element group 35: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_index_resize_1/index_resize_ack
      -- CP-element group 35: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_index_scale_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_index_scale_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_index_scale_1/scale_rename_req
      -- CP-element group 35: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_index_scale_1/scale_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_final_index_sum_regn_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_final_index_sum_regn_Sample/req
      -- 
    ca_6572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2609_inst_ack_1, ack => convTransposeD_CP_6285_elements(35)); -- 
    req_6597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(35), ack => array_obj_ref_2615_index_offset_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	55 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_final_index_sum_regn_sample_complete
      -- CP-element group 36: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_final_index_sum_regn_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_final_index_sum_regn_Sample/ack
      -- 
    ack_6598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2615_index_offset_ack_0, ack => convTransposeD_CP_6285_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	91 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (11) 
      -- CP-element group 37: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2616_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_offset_calculated
      -- CP-element group 37: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_final_index_sum_regn_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_final_index_sum_regn_Update/ack
      -- CP-element group 37: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_base_plus_offset/$entry
      -- CP-element group 37: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_base_plus_offset/$exit
      -- CP-element group 37: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_base_plus_offset/sum_rename_req
      -- CP-element group 37: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2616_request/$entry
      -- CP-element group 37: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2616_request/req
      -- 
    ack_6603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2615_index_offset_ack_1, ack => convTransposeD_CP_6285_elements(37)); -- 
    req_6612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(37), ack => addr_of_2616_final_reg_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2616_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2616_request/$exit
      -- CP-element group 38: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2616_request/ack
      -- 
    ack_6613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2616_final_reg_ack_0, ack => convTransposeD_CP_6285_elements(38)); -- 
    -- CP-element group 39:  join  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	91 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (24) 
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2616_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2616_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2616_complete/ack
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_base_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_word_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_base_address_resized
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_base_addr_resize/$entry
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_base_addr_resize/$exit
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_base_addr_resize/base_resize_req
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_base_addr_resize/base_resize_ack
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_word_addrgen/$entry
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_word_addrgen/$exit
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_word_addrgen/root_register_req
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_word_addrgen/root_register_ack
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_Sample/word_access_start/$entry
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_Sample/word_access_start/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_Sample/word_access_start/word_0/rr
      -- 
    ack_6618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2616_final_reg_ack_1, ack => convTransposeD_CP_6285_elements(39)); -- 
    rr_6651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(39), ack => ptr_deref_2620_load_0_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_Sample/word_access_start/$exit
      -- CP-element group 40: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_Sample/word_access_start/word_0/$exit
      -- CP-element group 40: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_Sample/word_access_start/word_0/ra
      -- 
    ra_6652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2620_load_0_ack_0, ack => convTransposeD_CP_6285_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	91 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	50 
    -- CP-element group 41:  members (9) 
      -- CP-element group 41: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_Update/word_access_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_Update/word_access_complete/word_0/$exit
      -- CP-element group 41: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_Update/word_access_complete/word_0/ca
      -- CP-element group 41: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_Update/ptr_deref_2620_Merge/$entry
      -- CP-element group 41: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_Update/ptr_deref_2620_Merge/$exit
      -- CP-element group 41: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_Update/ptr_deref_2620_Merge/merge_req
      -- CP-element group 41: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_Update/ptr_deref_2620_Merge/merge_ack
      -- 
    ca_6663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2620_load_0_ack_1, ack => convTransposeD_CP_6285_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	91 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2625_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2625_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2625_Sample/ra
      -- 
    ra_6677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2625_inst_ack_0, ack => convTransposeD_CP_6285_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	91 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2625_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2625_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2625_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2639_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2639_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2639_Sample/rr
      -- 
    ca_6682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2625_inst_ack_1, ack => convTransposeD_CP_6285_elements(43)); -- 
    rr_6690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(43), ack => type_cast_2639_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2639_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2639_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2639_Sample/ra
      -- 
    ra_6691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2639_inst_ack_0, ack => convTransposeD_CP_6285_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	91 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (16) 
      -- CP-element group 45: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_index_scale_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2639_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2639_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2639_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_index_resized_1
      -- CP-element group 45: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_index_scaled_1
      -- CP-element group 45: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_index_computed_1
      -- CP-element group 45: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_index_resize_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_index_resize_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_index_resize_1/index_resize_req
      -- CP-element group 45: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_index_resize_1/index_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_index_scale_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_index_scale_1/scale_rename_req
      -- CP-element group 45: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_index_scale_1/scale_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_final_index_sum_regn_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_final_index_sum_regn_Sample/req
      -- 
    ca_6696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2639_inst_ack_1, ack => convTransposeD_CP_6285_elements(45)); -- 
    req_6721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(45), ack => array_obj_ref_2645_index_offset_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	55 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_final_index_sum_regn_sample_complete
      -- CP-element group 46: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_final_index_sum_regn_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_final_index_sum_regn_Sample/ack
      -- 
    ack_6722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2645_index_offset_ack_0, ack => convTransposeD_CP_6285_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	91 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (11) 
      -- CP-element group 47: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2646_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_root_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_offset_calculated
      -- CP-element group 47: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_final_index_sum_regn_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_final_index_sum_regn_Update/ack
      -- CP-element group 47: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_base_plus_offset/$entry
      -- CP-element group 47: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_base_plus_offset/$exit
      -- CP-element group 47: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_base_plus_offset/sum_rename_req
      -- CP-element group 47: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_base_plus_offset/sum_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2646_request/$entry
      -- CP-element group 47: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2646_request/req
      -- 
    ack_6727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2645_index_offset_ack_1, ack => convTransposeD_CP_6285_elements(47)); -- 
    req_6736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(47), ack => addr_of_2646_final_reg_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2646_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2646_request/$exit
      -- CP-element group 48: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2646_request/ack
      -- 
    ack_6737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2646_final_reg_ack_0, ack => convTransposeD_CP_6285_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	91 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (19) 
      -- CP-element group 49: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2646_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2646_complete/$exit
      -- CP-element group 49: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2646_complete/ack
      -- CP-element group 49: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_base_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_word_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_base_address_resized
      -- CP-element group 49: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_base_addr_resize/$entry
      -- CP-element group 49: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_base_addr_resize/$exit
      -- CP-element group 49: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_base_addr_resize/base_resize_req
      -- CP-element group 49: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_base_addr_resize/base_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_word_addrgen/$entry
      -- CP-element group 49: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_word_addrgen/$exit
      -- CP-element group 49: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_word_addrgen/root_register_req
      -- CP-element group 49: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_word_addrgen/root_register_ack
      -- 
    ack_6742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2646_final_reg_ack_1, ack => convTransposeD_CP_6285_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	41 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_Sample/ptr_deref_2649_Split/$entry
      -- CP-element group 50: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_Sample/ptr_deref_2649_Split/$exit
      -- CP-element group 50: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_Sample/ptr_deref_2649_Split/split_req
      -- CP-element group 50: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_Sample/ptr_deref_2649_Split/split_ack
      -- CP-element group 50: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_Sample/word_access_start/$entry
      -- CP-element group 50: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_Sample/word_access_start/word_0/$entry
      -- CP-element group 50: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_Sample/word_access_start/word_0/rr
      -- 
    rr_6780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(50), ack => ptr_deref_2649_store_0_req_0); -- 
    convTransposeD_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6285_elements(41) & convTransposeD_CP_6285_elements(49);
      gj_convTransposeD_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6285_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_Sample/word_access_start/$exit
      -- CP-element group 51: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_Sample/word_access_start/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_Sample/word_access_start/word_0/ra
      -- 
    ra_6781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2649_store_0_ack_0, ack => convTransposeD_CP_6285_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	91 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_Update/word_access_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_Update/word_access_complete/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_Update/word_access_complete/word_0/ca
      -- 
    ca_6792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2649_store_0_ack_1, ack => convTransposeD_CP_6285_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	91 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2655_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2655_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2655_Sample/ra
      -- 
    ra_6801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2655_inst_ack_0, ack => convTransposeD_CP_6285_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	91 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2655_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2655_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2655_Update/ca
      -- 
    ca_6806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2655_inst_ack_1, ack => convTransposeD_CP_6285_elements(54)); -- 
    -- CP-element group 55:  branch  join  transition  place  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	52 
    -- CP-element group 55: 	54 
    -- CP-element group 55: 	36 
    -- CP-element group 55: 	46 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (10) 
      -- CP-element group 55: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669__exit__
      -- CP-element group 55: 	 branch_block_stmt_2417/if_stmt_2670__entry__
      -- CP-element group 55: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/$exit
      -- CP-element group 55: 	 branch_block_stmt_2417/if_stmt_2670_dead_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_2417/if_stmt_2670_eval_test/$entry
      -- CP-element group 55: 	 branch_block_stmt_2417/if_stmt_2670_eval_test/$exit
      -- CP-element group 55: 	 branch_block_stmt_2417/if_stmt_2670_eval_test/branch_req
      -- CP-element group 55: 	 branch_block_stmt_2417/R_cmp_2671_place
      -- CP-element group 55: 	 branch_block_stmt_2417/if_stmt_2670_if_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_2417/if_stmt_2670_else_link/$entry
      -- 
    branch_req_6814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(55), ack => if_stmt_2670_branch_req_0); -- 
    convTransposeD_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6285_elements(52) & convTransposeD_CP_6285_elements(54) & convTransposeD_CP_6285_elements(36) & convTransposeD_CP_6285_elements(46);
      gj_convTransposeD_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6285_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	86 
    -- CP-element group 56: 	87 
    -- CP-element group 56:  members (24) 
      -- CP-element group 56: 	 branch_block_stmt_2417/merge_stmt_2676__exit__
      -- CP-element group 56: 	 branch_block_stmt_2417/assign_stmt_2682__entry__
      -- CP-element group 56: 	 branch_block_stmt_2417/assign_stmt_2682__exit__
      -- CP-element group 56: 	 branch_block_stmt_2417/ifx_xthen_whilex_xbody
      -- CP-element group 56: 	 branch_block_stmt_2417/if_stmt_2670_if_link/$exit
      -- CP-element group 56: 	 branch_block_stmt_2417/if_stmt_2670_if_link/if_choice_transition
      -- CP-element group 56: 	 branch_block_stmt_2417/whilex_xbody_ifx_xthen
      -- CP-element group 56: 	 branch_block_stmt_2417/assign_stmt_2682/$entry
      -- CP-element group 56: 	 branch_block_stmt_2417/assign_stmt_2682/$exit
      -- CP-element group 56: 	 branch_block_stmt_2417/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_2417/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2568/$entry
      -- CP-element group 56: 	 branch_block_stmt_2417/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2568/phi_stmt_2568_sources/$entry
      -- CP-element group 56: 	 branch_block_stmt_2417/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2568/phi_stmt_2568_sources/type_cast_2571/$entry
      -- CP-element group 56: 	 branch_block_stmt_2417/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2568/phi_stmt_2568_sources/type_cast_2571/SplitProtocol/$entry
      -- CP-element group 56: 	 branch_block_stmt_2417/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2568/phi_stmt_2568_sources/type_cast_2571/SplitProtocol/Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_2417/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2568/phi_stmt_2568_sources/type_cast_2571/SplitProtocol/Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_2417/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2568/phi_stmt_2568_sources/type_cast_2571/SplitProtocol/Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_2417/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2568/phi_stmt_2568_sources/type_cast_2571/SplitProtocol/Update/cr
      -- CP-element group 56: 	 branch_block_stmt_2417/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_2417/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_2417/merge_stmt_2676_PhiReqMerge
      -- CP-element group 56: 	 branch_block_stmt_2417/merge_stmt_2676_PhiAck/$entry
      -- CP-element group 56: 	 branch_block_stmt_2417/merge_stmt_2676_PhiAck/$exit
      -- CP-element group 56: 	 branch_block_stmt_2417/merge_stmt_2676_PhiAck/dummy
      -- 
    if_choice_transition_6819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2670_branch_ack_1, ack => convTransposeD_CP_6285_elements(56)); -- 
    rr_7032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(56), ack => type_cast_2571_inst_req_0); -- 
    cr_7037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(56), ack => type_cast_2571_inst_req_1); -- 
    -- CP-element group 57:  fork  transition  place  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	59 
    -- CP-element group 57: 	61 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (24) 
      -- CP-element group 57: 	 branch_block_stmt_2417/merge_stmt_2684__exit__
      -- CP-element group 57: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725__entry__
      -- CP-element group 57: 	 branch_block_stmt_2417/if_stmt_2670_else_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_2417/if_stmt_2670_else_link/else_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_2417/whilex_xbody_ifx_xelse
      -- CP-element group 57: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/$entry
      -- CP-element group 57: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2694_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2694_update_start_
      -- CP-element group 57: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2694_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2694_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2694_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2694_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2709_update_start_
      -- CP-element group 57: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2709_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2709_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2719_update_start_
      -- CP-element group 57: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2719_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2719_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_2417/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_2417/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_2417/merge_stmt_2684_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_2417/merge_stmt_2684_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_2417/merge_stmt_2684_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_2417/merge_stmt_2684_PhiAck/dummy
      -- 
    else_choice_transition_6823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2670_branch_ack_0, ack => convTransposeD_CP_6285_elements(57)); -- 
    rr_6839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(57), ack => type_cast_2694_inst_req_0); -- 
    cr_6844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(57), ack => type_cast_2694_inst_req_1); -- 
    cr_6858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(57), ack => type_cast_2709_inst_req_1); -- 
    cr_6872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(57), ack => type_cast_2719_inst_req_1); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2694_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2694_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2694_Sample/ra
      -- 
    ra_6840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2694_inst_ack_0, ack => convTransposeD_CP_6285_elements(58)); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2694_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2694_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2694_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2709_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2709_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2709_Sample/rr
      -- 
    ca_6845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2694_inst_ack_1, ack => convTransposeD_CP_6285_elements(59)); -- 
    rr_6853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(59), ack => type_cast_2709_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2709_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2709_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2709_Sample/ra
      -- 
    ra_6854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2709_inst_ack_0, ack => convTransposeD_CP_6285_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	57 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2709_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2709_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2709_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2719_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2719_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2719_Sample/rr
      -- 
    ca_6859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2709_inst_ack_1, ack => convTransposeD_CP_6285_elements(61)); -- 
    rr_6867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(61), ack => type_cast_2719_inst_req_0); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2719_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2719_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2719_Sample/ra
      -- 
    ra_6868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2719_inst_ack_0, ack => convTransposeD_CP_6285_elements(62)); -- 
    -- CP-element group 63:  branch  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (13) 
      -- CP-element group 63: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725__exit__
      -- CP-element group 63: 	 branch_block_stmt_2417/if_stmt_2726__entry__
      -- CP-element group 63: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/$exit
      -- CP-element group 63: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2719_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2719_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_2417/assign_stmt_2690_to_assign_stmt_2725/type_cast_2719_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_2417/if_stmt_2726_dead_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_2417/if_stmt_2726_eval_test/$entry
      -- CP-element group 63: 	 branch_block_stmt_2417/if_stmt_2726_eval_test/$exit
      -- CP-element group 63: 	 branch_block_stmt_2417/if_stmt_2726_eval_test/branch_req
      -- CP-element group 63: 	 branch_block_stmt_2417/R_cmp137_2727_place
      -- CP-element group 63: 	 branch_block_stmt_2417/if_stmt_2726_if_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_2417/if_stmt_2726_else_link/$entry
      -- 
    ca_6873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2719_inst_ack_1, ack => convTransposeD_CP_6285_elements(63)); -- 
    branch_req_6881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(63), ack => if_stmt_2726_branch_req_0); -- 
    -- CP-element group 64:  merge  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (15) 
      -- CP-element group 64: 	 branch_block_stmt_2417/merge_stmt_2732__exit__
      -- CP-element group 64: 	 branch_block_stmt_2417/assign_stmt_2737__entry__
      -- CP-element group 64: 	 branch_block_stmt_2417/if_stmt_2726_if_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_2417/if_stmt_2726_if_link/if_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_2417/ifx_xelse_whilex_xend
      -- CP-element group 64: 	 branch_block_stmt_2417/assign_stmt_2737/$entry
      -- CP-element group 64: 	 branch_block_stmt_2417/assign_stmt_2737/WPIPE_Block3_done_2734_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_2417/assign_stmt_2737/WPIPE_Block3_done_2734_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_2417/assign_stmt_2737/WPIPE_Block3_done_2734_Sample/req
      -- CP-element group 64: 	 branch_block_stmt_2417/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_2417/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 64: 	 branch_block_stmt_2417/merge_stmt_2732_PhiReqMerge
      -- CP-element group 64: 	 branch_block_stmt_2417/merge_stmt_2732_PhiAck/$entry
      -- CP-element group 64: 	 branch_block_stmt_2417/merge_stmt_2732_PhiAck/$exit
      -- CP-element group 64: 	 branch_block_stmt_2417/merge_stmt_2732_PhiAck/dummy
      -- 
    if_choice_transition_6886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2726_branch_ack_1, ack => convTransposeD_CP_6285_elements(64)); -- 
    req_6903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(64), ack => WPIPE_Block3_done_2734_inst_req_0); -- 
    -- CP-element group 65:  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	75 
    -- CP-element group 65: 	76 
    -- CP-element group 65: 	78 
    -- CP-element group 65: 	79 
    -- CP-element group 65:  members (20) 
      -- CP-element group 65: 	 branch_block_stmt_2417/if_stmt_2726_else_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_2417/if_stmt_2726_else_link/else_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 65: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/$entry
      -- CP-element group 65: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/$entry
      -- CP-element group 65: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Update/cr
      -- CP-element group 65: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/$entry
      -- CP-element group 65: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/$entry
      -- CP-element group 65: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2726_branch_ack_0, ack => convTransposeD_CP_6285_elements(65)); -- 
    rr_6977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(65), ack => type_cast_2506_inst_req_0); -- 
    cr_6982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(65), ack => type_cast_2506_inst_req_1); -- 
    rr_7000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(65), ack => type_cast_2512_inst_req_0); -- 
    cr_7005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(65), ack => type_cast_2512_inst_req_1); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_2417/assign_stmt_2737/WPIPE_Block3_done_2734_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_2417/assign_stmt_2737/WPIPE_Block3_done_2734_update_start_
      -- CP-element group 66: 	 branch_block_stmt_2417/assign_stmt_2737/WPIPE_Block3_done_2734_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_2417/assign_stmt_2737/WPIPE_Block3_done_2734_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_2417/assign_stmt_2737/WPIPE_Block3_done_2734_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_2417/assign_stmt_2737/WPIPE_Block3_done_2734_Update/req
      -- 
    ack_6904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2734_inst_ack_0, ack => convTransposeD_CP_6285_elements(66)); -- 
    req_6908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(66), ack => WPIPE_Block3_done_2734_inst_req_1); -- 
    -- CP-element group 67:  transition  place  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (16) 
      -- CP-element group 67: 	 $exit
      -- CP-element group 67: 	 branch_block_stmt_2417/$exit
      -- CP-element group 67: 	 branch_block_stmt_2417/branch_block_stmt_2417__exit__
      -- CP-element group 67: 	 branch_block_stmt_2417/assign_stmt_2737__exit__
      -- CP-element group 67: 	 branch_block_stmt_2417/return__
      -- CP-element group 67: 	 branch_block_stmt_2417/merge_stmt_2739__exit__
      -- CP-element group 67: 	 branch_block_stmt_2417/assign_stmt_2737/$exit
      -- CP-element group 67: 	 branch_block_stmt_2417/assign_stmt_2737/WPIPE_Block3_done_2734_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_2417/assign_stmt_2737/WPIPE_Block3_done_2734_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_2417/assign_stmt_2737/WPIPE_Block3_done_2734_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_2417/return___PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2417/return___PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_2417/merge_stmt_2739_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_2417/merge_stmt_2739_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_2417/merge_stmt_2739_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_2417/merge_stmt_2739_PhiAck/dummy
      -- 
    ack_6909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2734_inst_ack_1, ack => convTransposeD_CP_6285_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	31 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Sample/ra
      -- 
    ra_6929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2508_inst_ack_0, ack => convTransposeD_CP_6285_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	31 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Update/ca
      -- 
    ca_6934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2508_inst_ack_1, ack => convTransposeD_CP_6285_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (5) 
      -- CP-element group 70: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/$exit
      -- CP-element group 70: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/$exit
      -- CP-element group 70: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/$exit
      -- CP-element group 70: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/$exit
      -- CP-element group 70: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_req
      -- 
    phi_stmt_2503_req_6935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2503_req_6935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(70), ack => phi_stmt_2503_req_1); -- 
    convTransposeD_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6285_elements(68) & convTransposeD_CP_6285_elements(69);
      gj_convTransposeD_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6285_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	31 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2514/SplitProtocol/Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2514/SplitProtocol/Sample/ra
      -- 
    ra_6952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2514_inst_ack_0, ack => convTransposeD_CP_6285_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	31 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2514/SplitProtocol/Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2514/SplitProtocol/Update/ca
      -- 
    ca_6957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2514_inst_ack_1, ack => convTransposeD_CP_6285_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/$exit
      -- CP-element group 73: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/$exit
      -- CP-element group 73: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2514/$exit
      -- CP-element group 73: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2514/SplitProtocol/$exit
      -- CP-element group 73: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_req
      -- 
    phi_stmt_2509_req_6958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2509_req_6958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(73), ack => phi_stmt_2509_req_1); -- 
    convTransposeD_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6285_elements(71) & convTransposeD_CP_6285_elements(72);
      gj_convTransposeD_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6285_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	82 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_2417/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6285_elements(70) & convTransposeD_CP_6285_elements(73);
      gj_convTransposeD_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6285_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	65 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Sample/ra
      -- 
    ra_6978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2506_inst_ack_0, ack => convTransposeD_CP_6285_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	65 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Update/ca
      -- 
    ca_6983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2506_inst_ack_1, ack => convTransposeD_CP_6285_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	81 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/$exit
      -- CP-element group 77: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/$exit
      -- CP-element group 77: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/$exit
      -- CP-element group 77: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2503/phi_stmt_2503_req
      -- 
    phi_stmt_2503_req_6984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2503_req_6984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(77), ack => phi_stmt_2503_req_0); -- 
    convTransposeD_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6285_elements(75) & convTransposeD_CP_6285_elements(76);
      gj_convTransposeD_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6285_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	65 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Sample/ra
      -- 
    ra_7001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2512_inst_ack_0, ack => convTransposeD_CP_6285_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	65 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/Update/ca
      -- 
    ca_7006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2512_inst_ack_1, ack => convTransposeD_CP_6285_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/$exit
      -- CP-element group 80: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/$exit
      -- CP-element group 80: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2512/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2509/phi_stmt_2509_req
      -- 
    phi_stmt_2509_req_7007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2509_req_7007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(80), ack => phi_stmt_2509_req_0); -- 
    convTransposeD_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6285_elements(78) & convTransposeD_CP_6285_elements(79);
      gj_convTransposeD_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6285_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	77 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2417/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6285_elements(77) & convTransposeD_CP_6285_elements(80);
      gj_convTransposeD_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6285_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  merge  fork  transition  place  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	74 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2417/merge_stmt_2502_PhiReqMerge
      -- CP-element group 82: 	 branch_block_stmt_2417/merge_stmt_2502_PhiAck/$entry
      -- 
    convTransposeD_CP_6285_elements(82) <= OrReduce(convTransposeD_CP_6285_elements(74) & convTransposeD_CP_6285_elements(81));
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_2417/merge_stmt_2502_PhiAck/phi_stmt_2503_ack
      -- 
    phi_stmt_2503_ack_7012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2503_ack_0, ack => convTransposeD_CP_6285_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_2417/merge_stmt_2502_PhiAck/phi_stmt_2509_ack
      -- 
    phi_stmt_2509_ack_7013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2509_ack_0, ack => convTransposeD_CP_6285_elements(84)); -- 
    -- CP-element group 85:  join  transition  place  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	89 
    -- CP-element group 85:  members (10) 
      -- CP-element group 85: 	 branch_block_stmt_2417/merge_stmt_2502__exit__
      -- CP-element group 85: 	 branch_block_stmt_2417/assign_stmt_2520_to_assign_stmt_2565__entry__
      -- CP-element group 85: 	 branch_block_stmt_2417/assign_stmt_2520_to_assign_stmt_2565__exit__
      -- CP-element group 85: 	 branch_block_stmt_2417/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 85: 	 branch_block_stmt_2417/assign_stmt_2520_to_assign_stmt_2565/$entry
      -- CP-element group 85: 	 branch_block_stmt_2417/assign_stmt_2520_to_assign_stmt_2565/$exit
      -- CP-element group 85: 	 branch_block_stmt_2417/merge_stmt_2502_PhiAck/$exit
      -- CP-element group 85: 	 branch_block_stmt_2417/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 85: 	 branch_block_stmt_2417/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2568/$entry
      -- CP-element group 85: 	 branch_block_stmt_2417/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2568/phi_stmt_2568_sources/$entry
      -- 
    convTransposeD_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6285_elements(83) & convTransposeD_CP_6285_elements(84);
      gj_convTransposeD_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6285_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	56 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2417/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2568/phi_stmt_2568_sources/type_cast_2571/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_2417/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2568/phi_stmt_2568_sources/type_cast_2571/SplitProtocol/Sample/ra
      -- 
    ra_7033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2571_inst_ack_0, ack => convTransposeD_CP_6285_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	56 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_2417/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2568/phi_stmt_2568_sources/type_cast_2571/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_2417/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2568/phi_stmt_2568_sources/type_cast_2571/SplitProtocol/Update/ca
      -- 
    ca_7038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2571_inst_ack_1, ack => convTransposeD_CP_6285_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (6) 
      -- CP-element group 88: 	 branch_block_stmt_2417/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 88: 	 branch_block_stmt_2417/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2568/$exit
      -- CP-element group 88: 	 branch_block_stmt_2417/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2568/phi_stmt_2568_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_2417/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2568/phi_stmt_2568_sources/type_cast_2571/$exit
      -- CP-element group 88: 	 branch_block_stmt_2417/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2568/phi_stmt_2568_sources/type_cast_2571/SplitProtocol/$exit
      -- CP-element group 88: 	 branch_block_stmt_2417/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2568/phi_stmt_2568_req
      -- 
    phi_stmt_2568_req_7039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2568_req_7039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(88), ack => phi_stmt_2568_req_0); -- 
    convTransposeD_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6285_elements(86) & convTransposeD_CP_6285_elements(87);
      gj_convTransposeD_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6285_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  output  delay-element  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	85 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_2417/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 89: 	 branch_block_stmt_2417/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2568/$exit
      -- CP-element group 89: 	 branch_block_stmt_2417/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2568/phi_stmt_2568_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_2417/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2568/phi_stmt_2568_sources/type_cast_2574_konst_delay_trans
      -- CP-element group 89: 	 branch_block_stmt_2417/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2568/phi_stmt_2568_req
      -- 
    phi_stmt_2568_req_7050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2568_req_7050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(89), ack => phi_stmt_2568_req_1); -- 
    -- Element group convTransposeD_CP_6285_elements(89) is a control-delay.
    cp_element_89_delay: control_delay_element  generic map(name => " 89_delay", delay_value => 1)  port map(req => convTransposeD_CP_6285_elements(85), ack => convTransposeD_CP_6285_elements(89), clk => clk, reset =>reset);
    -- CP-element group 90:  merge  transition  place  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_2417/merge_stmt_2567_PhiReqMerge
      -- CP-element group 90: 	 branch_block_stmt_2417/merge_stmt_2567_PhiAck/$entry
      -- 
    convTransposeD_CP_6285_elements(90) <= OrReduce(convTransposeD_CP_6285_elements(88) & convTransposeD_CP_6285_elements(89));
    -- CP-element group 91:  fork  transition  place  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	52 
    -- CP-element group 91: 	53 
    -- CP-element group 91: 	54 
    -- CP-element group 91: 	41 
    -- CP-element group 91: 	42 
    -- CP-element group 91: 	43 
    -- CP-element group 91: 	45 
    -- CP-element group 91: 	32 
    -- CP-element group 91: 	33 
    -- CP-element group 91: 	35 
    -- CP-element group 91: 	37 
    -- CP-element group 91: 	39 
    -- CP-element group 91: 	47 
    -- CP-element group 91: 	49 
    -- CP-element group 91:  members (51) 
      -- CP-element group 91: 	 branch_block_stmt_2417/merge_stmt_2567__exit__
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669__entry__
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/$entry
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2595_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2595_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2595_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2595_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2595_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2595_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2609_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2609_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2609_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2616_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_final_index_sum_regn_update_start
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_final_index_sum_regn_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2615_final_index_sum_regn_Update/req
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2616_complete/$entry
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2616_complete/req
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_Update/word_access_complete/$entry
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_Update/word_access_complete/word_0/$entry
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2620_Update/word_access_complete/word_0/cr
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2625_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2625_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2625_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2625_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2625_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2625_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2639_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2639_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2639_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2646_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_final_index_sum_regn_update_start
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_final_index_sum_regn_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/array_obj_ref_2645_final_index_sum_regn_Update/req
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2646_complete/$entry
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/addr_of_2646_complete/req
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_Update/word_access_complete/$entry
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_Update/word_access_complete/word_0/$entry
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/ptr_deref_2649_Update/word_access_complete/word_0/cr
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2655_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2655_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2655_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2655_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2655_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2417/assign_stmt_2581_to_assign_stmt_2669/type_cast_2655_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_2417/merge_stmt_2567_PhiAck/$exit
      -- CP-element group 91: 	 branch_block_stmt_2417/merge_stmt_2567_PhiAck/phi_stmt_2568_ack
      -- 
    phi_stmt_2568_ack_7055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2568_ack_0, ack => convTransposeD_CP_6285_elements(91)); -- 
    rr_6552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(91), ack => type_cast_2595_inst_req_0); -- 
    cr_6557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(91), ack => type_cast_2595_inst_req_1); -- 
    cr_6571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(91), ack => type_cast_2609_inst_req_1); -- 
    req_6602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(91), ack => array_obj_ref_2615_index_offset_req_1); -- 
    req_6617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(91), ack => addr_of_2616_final_reg_req_1); -- 
    cr_6662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(91), ack => ptr_deref_2620_load_0_req_1); -- 
    rr_6676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(91), ack => type_cast_2625_inst_req_0); -- 
    cr_6681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(91), ack => type_cast_2625_inst_req_1); -- 
    cr_6695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(91), ack => type_cast_2639_inst_req_1); -- 
    req_6726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(91), ack => array_obj_ref_2645_index_offset_req_1); -- 
    req_6741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(91), ack => addr_of_2646_final_reg_req_1); -- 
    cr_6791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(91), ack => ptr_deref_2649_store_0_req_1); -- 
    rr_6800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(91), ack => type_cast_2655_inst_req_0); -- 
    cr_6805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6285_elements(91), ack => type_cast_2655_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2603_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2633_wire : std_logic_vector(31 downto 0);
    signal R_idxprom102_2644_resized : std_logic_vector(13 downto 0);
    signal R_idxprom102_2644_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2614_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2614_scaled : std_logic_vector(13 downto 0);
    signal add107_2662 : std_logic_vector(31 downto 0);
    signal add49_2586 : std_logic_vector(15 downto 0);
    signal add93_2591 : std_logic_vector(15 downto 0);
    signal array_obj_ref_2615_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2615_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2615_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2615_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2615_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2615_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2645_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2645_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2645_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2645_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2645_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2645_root_address : std_logic_vector(13 downto 0);
    signal arrayidx103_2647 : std_logic_vector(31 downto 0);
    signal arrayidx97_2617 : std_logic_vector(31 downto 0);
    signal call11_2438 : std_logic_vector(15 downto 0);
    signal call13_2441 : std_logic_vector(15 downto 0);
    signal call14_2444 : std_logic_vector(15 downto 0);
    signal call15_2447 : std_logic_vector(15 downto 0);
    signal call17_2450 : std_logic_vector(15 downto 0);
    signal call19_2453 : std_logic_vector(15 downto 0);
    signal call1_2423 : std_logic_vector(15 downto 0);
    signal call3_2426 : std_logic_vector(15 downto 0);
    signal call5_2429 : std_logic_vector(15 downto 0);
    signal call7_2432 : std_logic_vector(15 downto 0);
    signal call9_2435 : std_logic_vector(15 downto 0);
    signal call_2420 : std_logic_vector(15 downto 0);
    signal cmp122_2700 : std_logic_vector(0 downto 0);
    signal cmp137_2725 : std_logic_vector(0 downto 0);
    signal cmp_2669 : std_logic_vector(0 downto 0);
    signal conv100_2626 : std_logic_vector(31 downto 0);
    signal conv106_2656 : std_logic_vector(31 downto 0);
    signal conv110_2470 : std_logic_vector(31 downto 0);
    signal conv118_2695 : std_logic_vector(31 downto 0);
    signal conv121_2474 : std_logic_vector(31 downto 0);
    signal conv133_2720 : std_logic_vector(31 downto 0);
    signal conv136_2478 : std_logic_vector(31 downto 0);
    signal conv96_2596 : std_logic_vector(31 downto 0);
    signal div27_2466 : std_logic_vector(15 downto 0);
    signal div_2460 : std_logic_vector(15 downto 0);
    signal idxprom102_2640 : std_logic_vector(63 downto 0);
    signal idxprom_2610 : std_logic_vector(63 downto 0);
    signal inc126_2710 : std_logic_vector(15 downto 0);
    signal inc_2690 : std_logic_vector(15 downto 0);
    signal indvar_2568 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2682 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_2715 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2509 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2503 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2706 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2581 : std_logic_vector(15 downto 0);
    signal ptr_deref_2620_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2620_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2620_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2620_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2620_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2649_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2649_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2649_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2649_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2649_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2649_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr101_2635 : std_logic_vector(31 downto 0);
    signal shr_2605 : std_logic_vector(31 downto 0);
    signal tmp10_2565 : std_logic_vector(15 downto 0);
    signal tmp164_2520 : std_logic_vector(15 downto 0);
    signal tmp165_2525 : std_logic_vector(15 downto 0);
    signal tmp166_2530 : std_logic_vector(15 downto 0);
    signal tmp1_2489 : std_logic_vector(15 downto 0);
    signal tmp2_2535 : std_logic_vector(15 downto 0);
    signal tmp3_2540 : std_logic_vector(15 downto 0);
    signal tmp4_2495 : std_logic_vector(15 downto 0);
    signal tmp5_2500 : std_logic_vector(15 downto 0);
    signal tmp6_2545 : std_logic_vector(15 downto 0);
    signal tmp7_2550 : std_logic_vector(15 downto 0);
    signal tmp8_2555 : std_logic_vector(15 downto 0);
    signal tmp98_2621 : std_logic_vector(63 downto 0);
    signal tmp9_2560 : std_logic_vector(15 downto 0);
    signal tmp_2484 : std_logic_vector(15 downto 0);
    signal type_cast_2458_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2464_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2482_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2493_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2506_wire : std_logic_vector(15 downto 0);
    signal type_cast_2508_wire : std_logic_vector(15 downto 0);
    signal type_cast_2512_wire : std_logic_vector(15 downto 0);
    signal type_cast_2514_wire : std_logic_vector(15 downto 0);
    signal type_cast_2571_wire : std_logic_vector(15 downto 0);
    signal type_cast_2574_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2579_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2594_wire : std_logic_vector(31 downto 0);
    signal type_cast_2599_wire : std_logic_vector(31 downto 0);
    signal type_cast_2602_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2608_wire : std_logic_vector(63 downto 0);
    signal type_cast_2624_wire : std_logic_vector(31 downto 0);
    signal type_cast_2629_wire : std_logic_vector(31 downto 0);
    signal type_cast_2632_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2638_wire : std_logic_vector(63 downto 0);
    signal type_cast_2654_wire : std_logic_vector(31 downto 0);
    signal type_cast_2660_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2665_wire : std_logic_vector(31 downto 0);
    signal type_cast_2667_wire : std_logic_vector(31 downto 0);
    signal type_cast_2680_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2688_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2693_wire : std_logic_vector(31 downto 0);
    signal type_cast_2718_wire : std_logic_vector(31 downto 0);
    signal type_cast_2736_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2615_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2615_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2615_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2615_resized_base_address <= "00000000000000";
    array_obj_ref_2645_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2645_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2645_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2645_resized_base_address <= "00000000000000";
    ptr_deref_2620_word_offset_0 <= "00000000000000";
    ptr_deref_2649_word_offset_0 <= "00000000000000";
    type_cast_2458_wire_constant <= "0000000000000001";
    type_cast_2464_wire_constant <= "0000000000000001";
    type_cast_2482_wire_constant <= "1111111111111111";
    type_cast_2493_wire_constant <= "1111111111111111";
    type_cast_2574_wire_constant <= "0000000000000000";
    type_cast_2579_wire_constant <= "0000000000000100";
    type_cast_2602_wire_constant <= "00000000000000000000000000000010";
    type_cast_2632_wire_constant <= "00000000000000000000000000000010";
    type_cast_2660_wire_constant <= "00000000000000000000000000000100";
    type_cast_2680_wire_constant <= "0000000000000001";
    type_cast_2688_wire_constant <= "0000000000000001";
    type_cast_2736_wire_constant <= "0000000000000001";
    phi_stmt_2503: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2506_wire & type_cast_2508_wire;
      req <= phi_stmt_2503_req_0 & phi_stmt_2503_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2503",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2503_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2503,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2503
    phi_stmt_2509: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2512_wire & type_cast_2514_wire;
      req <= phi_stmt_2509_req_0 & phi_stmt_2509_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2509",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2509_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2509,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2509
    phi_stmt_2568: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2571_wire & type_cast_2574_wire_constant;
      req <= phi_stmt_2568_req_0 & phi_stmt_2568_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2568",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2568_ack_0,
          idata => idata,
          odata => indvar_2568,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2568
    -- flow-through select operator MUX_2705_inst
    input_dim1x_x2_2706 <= div27_2466 when (cmp122_2700(0) /=  '0') else inc_2690;
    addr_of_2616_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2616_final_reg_req_0;
      addr_of_2616_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2616_final_reg_req_1;
      addr_of_2616_final_reg_ack_1<= rack(0);
      addr_of_2616_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2616_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2615_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx97_2617,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2646_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2646_final_reg_req_0;
      addr_of_2646_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2646_final_reg_req_1;
      addr_of_2646_final_reg_ack_1<= rack(0);
      addr_of_2646_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2646_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2645_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx103_2647,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2469_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2469_inst_req_0;
      type_cast_2469_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2469_inst_req_1;
      type_cast_2469_inst_ack_1<= rack(0);
      type_cast_2469_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2469_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2426,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv110_2470,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2473_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2473_inst_req_0;
      type_cast_2473_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2473_inst_req_1;
      type_cast_2473_inst_ack_1<= rack(0);
      type_cast_2473_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2473_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_2423,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv121_2474,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2477_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2477_inst_req_0;
      type_cast_2477_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2477_inst_req_1;
      type_cast_2477_inst_ack_1<= rack(0);
      type_cast_2477_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2477_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2420,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv136_2478,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2506_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2506_inst_req_0;
      type_cast_2506_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2506_inst_req_1;
      type_cast_2506_inst_ack_1<= rack(0);
      type_cast_2506_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2506_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2706,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2506_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2508_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2508_inst_req_0;
      type_cast_2508_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2508_inst_req_1;
      type_cast_2508_inst_ack_1<= rack(0);
      type_cast_2508_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2508_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div27_2466,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2508_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2512_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2512_inst_req_0;
      type_cast_2512_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2512_inst_req_1;
      type_cast_2512_inst_ack_1<= rack(0);
      type_cast_2512_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2512_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_2715,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2512_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2514_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2514_inst_req_0;
      type_cast_2514_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2514_inst_req_1;
      type_cast_2514_inst_ack_1<= rack(0);
      type_cast_2514_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2514_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2460,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2514_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2571_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2571_inst_req_0;
      type_cast_2571_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2571_inst_req_1;
      type_cast_2571_inst_ack_1<= rack(0);
      type_cast_2571_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2571_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2682,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2571_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2595_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2595_inst_req_0;
      type_cast_2595_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2595_inst_req_1;
      type_cast_2595_inst_ack_1<= rack(0);
      type_cast_2595_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2595_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2594_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv96_2596,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2599_inst
    process(conv96_2596) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv96_2596(31 downto 0);
      type_cast_2599_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2604_inst
    process(ASHR_i32_i32_2603_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2603_wire(31 downto 0);
      shr_2605 <= tmp_var; -- 
    end process;
    type_cast_2609_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2609_inst_req_0;
      type_cast_2609_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2609_inst_req_1;
      type_cast_2609_inst_ack_1<= rack(0);
      type_cast_2609_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2609_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2608_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2610,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2625_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2625_inst_req_0;
      type_cast_2625_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2625_inst_req_1;
      type_cast_2625_inst_ack_1<= rack(0);
      type_cast_2625_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2625_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2624_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv100_2626,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2629_inst
    process(conv100_2626) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv100_2626(31 downto 0);
      type_cast_2629_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2634_inst
    process(ASHR_i32_i32_2633_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2633_wire(31 downto 0);
      shr101_2635 <= tmp_var; -- 
    end process;
    type_cast_2639_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2639_inst_req_0;
      type_cast_2639_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2639_inst_req_1;
      type_cast_2639_inst_ack_1<= rack(0);
      type_cast_2639_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2639_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2638_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom102_2640,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2655_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2655_inst_req_0;
      type_cast_2655_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2655_inst_req_1;
      type_cast_2655_inst_ack_1<= rack(0);
      type_cast_2655_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2655_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2654_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv106_2656,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2665_inst
    process(add107_2662) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add107_2662(31 downto 0);
      type_cast_2665_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2667_inst
    process(conv110_2470) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv110_2470(31 downto 0);
      type_cast_2667_wire <= tmp_var; -- 
    end process;
    type_cast_2694_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2694_inst_req_0;
      type_cast_2694_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2694_inst_req_1;
      type_cast_2694_inst_ack_1<= rack(0);
      type_cast_2694_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2694_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2693_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv118_2695,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2709_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2709_inst_req_0;
      type_cast_2709_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2709_inst_req_1;
      type_cast_2709_inst_ack_1<= rack(0);
      type_cast_2709_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2709_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp122_2700,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc126_2710,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2719_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2719_inst_req_0;
      type_cast_2719_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2719_inst_req_1;
      type_cast_2719_inst_ack_1<= rack(0);
      type_cast_2719_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2719_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2718_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv133_2720,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2615_index_1_rename
    process(R_idxprom_2614_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2614_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2614_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2615_index_1_resize
    process(idxprom_2610) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2610;
      ov := iv(13 downto 0);
      R_idxprom_2614_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2615_root_address_inst
    process(array_obj_ref_2615_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2615_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2615_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2645_index_1_rename
    process(R_idxprom102_2644_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom102_2644_resized;
      ov(13 downto 0) := iv;
      R_idxprom102_2644_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2645_index_1_resize
    process(idxprom102_2640) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom102_2640;
      ov := iv(13 downto 0);
      R_idxprom102_2644_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2645_root_address_inst
    process(array_obj_ref_2645_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2645_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2645_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2620_addr_0
    process(ptr_deref_2620_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2620_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2620_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2620_base_resize
    process(arrayidx97_2617) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx97_2617;
      ov := iv(13 downto 0);
      ptr_deref_2620_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2620_gather_scatter
    process(ptr_deref_2620_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2620_data_0;
      ov(63 downto 0) := iv;
      tmp98_2621 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2620_root_address_inst
    process(ptr_deref_2620_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2620_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2620_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2649_addr_0
    process(ptr_deref_2649_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2649_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2649_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2649_base_resize
    process(arrayidx103_2647) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx103_2647;
      ov := iv(13 downto 0);
      ptr_deref_2649_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2649_gather_scatter
    process(tmp98_2621) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp98_2621;
      ov(63 downto 0) := iv;
      ptr_deref_2649_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2649_root_address_inst
    process(ptr_deref_2649_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2649_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2649_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2670_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2669;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2670_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2670_branch_req_0,
          ack0 => if_stmt_2670_branch_ack_0,
          ack1 => if_stmt_2670_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2726_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp137_2725;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2726_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2726_branch_req_0,
          ack0 => if_stmt_2726_branch_ack_0,
          ack1 => if_stmt_2726_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2483_inst
    process(call9_2435) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2435, type_cast_2482_wire_constant, tmp_var);
      tmp_2484 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2494_inst
    process(call7_2432) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2432, type_cast_2493_wire_constant, tmp_var);
      tmp4_2495 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2524_inst
    process(input_dim1x_x1x_xph_2503, tmp164_2520) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2503, tmp164_2520, tmp_var);
      tmp165_2525 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2539_inst
    process(tmp1_2489, tmp2_2535) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp1_2489, tmp2_2535, tmp_var);
      tmp3_2540 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2549_inst
    process(tmp5_2500, tmp6_2545) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp5_2500, tmp6_2545, tmp_var);
      tmp7_2550 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2559_inst
    process(tmp3_2540, tmp8_2555) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_2540, tmp8_2555, tmp_var);
      tmp9_2560 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2585_inst
    process(tmp166_2530, input_dim2x_x1_2581) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp166_2530, input_dim2x_x1_2581, tmp_var);
      add49_2586 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2590_inst
    process(tmp10_2565, input_dim2x_x1_2581) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp10_2565, input_dim2x_x1_2581, tmp_var);
      add93_2591 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2681_inst
    process(indvar_2568) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2568, type_cast_2680_wire_constant, tmp_var);
      indvarx_xnext_2682 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2689_inst
    process(input_dim1x_x1x_xph_2503) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2503, type_cast_2688_wire_constant, tmp_var);
      inc_2690 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2714_inst
    process(inc126_2710, input_dim0x_x2x_xph_2509) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc126_2710, input_dim0x_x2x_xph_2509, tmp_var);
      input_dim0x_x0_2715 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2661_inst
    process(conv106_2656) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv106_2656, type_cast_2660_wire_constant, tmp_var);
      add107_2662 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2603_inst
    process(type_cast_2599_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2599_wire, type_cast_2602_wire_constant, tmp_var);
      ASHR_i32_i32_2603_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2633_inst
    process(type_cast_2629_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2629_wire, type_cast_2632_wire_constant, tmp_var);
      ASHR_i32_i32_2633_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2699_inst
    process(conv118_2695, conv121_2474) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv118_2695, conv121_2474, tmp_var);
      cmp122_2700 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2724_inst
    process(conv133_2720, conv136_2478) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv133_2720, conv136_2478, tmp_var);
      cmp137_2725 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2459_inst
    process(call_2420) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2420, type_cast_2458_wire_constant, tmp_var);
      div_2460 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2465_inst
    process(call1_2423) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call1_2423, type_cast_2464_wire_constant, tmp_var);
      div27_2466 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2519_inst
    process(call1_2423, input_dim0x_x2x_xph_2509) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call1_2423, input_dim0x_x2x_xph_2509, tmp_var);
      tmp164_2520 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2529_inst
    process(call3_2426, tmp165_2525) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call3_2426, tmp165_2525, tmp_var);
      tmp166_2530 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2534_inst
    process(call13_2441, input_dim1x_x1x_xph_2503) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_2441, input_dim1x_x1x_xph_2503, tmp_var);
      tmp2_2535 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2544_inst
    process(call13_2441, input_dim0x_x2x_xph_2509) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_2441, input_dim0x_x2x_xph_2509, tmp_var);
      tmp6_2545 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2554_inst
    process(call17_2450, tmp7_2550) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call17_2450, tmp7_2550, tmp_var);
      tmp8_2555 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2564_inst
    process(call19_2453, tmp9_2560) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call19_2453, tmp9_2560, tmp_var);
      tmp10_2565 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2580_inst
    process(indvar_2568) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2568, type_cast_2579_wire_constant, tmp_var);
      input_dim2x_x1_2581 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2668_inst
    process(type_cast_2665_wire, type_cast_2667_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2665_wire, type_cast_2667_wire, tmp_var);
      cmp_2669 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2488_inst
    process(tmp_2484, call14_2444) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp_2484, call14_2444, tmp_var);
      tmp1_2489 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2499_inst
    process(tmp4_2495, call14_2444) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp4_2495, call14_2444, tmp_var);
      tmp5_2500 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_2615_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2614_scaled;
      array_obj_ref_2615_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2615_index_offset_req_0;
      array_obj_ref_2615_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2615_index_offset_req_1;
      array_obj_ref_2615_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_2645_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom102_2644_scaled;
      array_obj_ref_2645_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2645_index_offset_req_0;
      array_obj_ref_2645_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2645_index_offset_req_1;
      array_obj_ref_2645_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- unary operator type_cast_2594_inst
    process(add49_2586) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add49_2586, tmp_var);
      type_cast_2594_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2608_inst
    process(shr_2605) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2605, tmp_var);
      type_cast_2608_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2624_inst
    process(add93_2591) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add93_2591, tmp_var);
      type_cast_2624_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2638_inst
    process(shr101_2635) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr101_2635, tmp_var);
      type_cast_2638_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2654_inst
    process(input_dim2x_x1_2581) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_2581, tmp_var);
      type_cast_2654_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2693_inst
    process(inc_2690) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2690, tmp_var);
      type_cast_2693_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2718_inst
    process(input_dim0x_x0_2715) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x0_2715, tmp_var);
      type_cast_2718_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_2620_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2620_load_0_req_0;
      ptr_deref_2620_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2620_load_0_req_1;
      ptr_deref_2620_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2620_word_address_0;
      ptr_deref_2620_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2649_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2649_store_0_req_0;
      ptr_deref_2649_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2649_store_0_req_1;
      ptr_deref_2649_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2649_word_address_0;
      data_in <= ptr_deref_2649_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_start_2440_inst RPIPE_Block3_start_2443_inst RPIPE_Block3_start_2446_inst RPIPE_Block3_start_2449_inst RPIPE_Block3_start_2452_inst RPIPE_Block3_start_2437_inst RPIPE_Block3_start_2434_inst RPIPE_Block3_start_2431_inst RPIPE_Block3_start_2428_inst RPIPE_Block3_start_2425_inst RPIPE_Block3_start_2422_inst RPIPE_Block3_start_2419_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(191 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 11 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 11 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant outBUFs : IntegerArray(11 downto 0) := (11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      reqL_unguarded(11) <= RPIPE_Block3_start_2440_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block3_start_2443_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block3_start_2446_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block3_start_2449_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block3_start_2452_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block3_start_2437_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block3_start_2434_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block3_start_2431_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block3_start_2428_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block3_start_2425_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block3_start_2422_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block3_start_2419_inst_req_0;
      RPIPE_Block3_start_2440_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block3_start_2443_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block3_start_2446_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block3_start_2449_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block3_start_2452_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block3_start_2437_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block3_start_2434_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block3_start_2431_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block3_start_2428_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block3_start_2425_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block3_start_2422_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block3_start_2419_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(11) <= RPIPE_Block3_start_2440_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block3_start_2443_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block3_start_2446_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block3_start_2449_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block3_start_2452_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block3_start_2437_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block3_start_2434_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block3_start_2431_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block3_start_2428_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block3_start_2425_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block3_start_2422_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block3_start_2419_inst_req_1;
      RPIPE_Block3_start_2440_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block3_start_2443_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block3_start_2446_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block3_start_2449_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block3_start_2452_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block3_start_2437_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block3_start_2434_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block3_start_2431_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block3_start_2428_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block3_start_2425_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block3_start_2422_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block3_start_2419_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      call13_2441 <= data_out(191 downto 176);
      call14_2444 <= data_out(175 downto 160);
      call15_2447 <= data_out(159 downto 144);
      call17_2450 <= data_out(143 downto 128);
      call19_2453 <= data_out(127 downto 112);
      call11_2438 <= data_out(111 downto 96);
      call9_2435 <= data_out(95 downto 80);
      call7_2432 <= data_out(79 downto 64);
      call5_2429 <= data_out(63 downto 48);
      call3_2426 <= data_out(47 downto 32);
      call1_2423 <= data_out(31 downto 16);
      call_2420 <= data_out(15 downto 0);
      Block3_start_read_0_gI: SplitGuardInterface generic map(name => "Block3_start_read_0_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_start_read_0: InputPortRevised -- 
        generic map ( name => "Block3_start_read_0", data_width => 16,  num_reqs => 12,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_start_pipe_read_req(0),
          oack => Block3_start_pipe_read_ack(0),
          odata => Block3_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_2734_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_2734_inst_req_0;
      WPIPE_Block3_done_2734_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_2734_inst_req_1;
      WPIPE_Block3_done_2734_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2736_wire_constant;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_29_load_0_req_0 : boolean;
  signal LOAD_count_29_load_0_ack_0 : boolean;
  signal LOAD_count_29_load_0_req_1 : boolean;
  signal LOAD_count_29_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Update/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_30/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_sample_start_
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_update_start_
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Sample/$entry
      -- 
    rr_21_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_21_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_29_load_0_req_0); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_29_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_sample_completed_
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_Sample/$exit
      -- 
    ra_22_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_29_load_0_ack_0, ack => timer_CP_0_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/LOAD_count_29_Merge/$entry
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_30/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_update_completed_
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/LOAD_count_29_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/LOAD_count_29_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/LOAD_count_29_Merge/merge_ack
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_29_load_0_ack_1, ack => timer_CP_0_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_29_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_29_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_29_word_address_0 <= "0";
    -- equivalence LOAD_count_29_gather_scatter
    process(LOAD_count_29_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_29_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_29_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_29_load_0_req_0;
      LOAD_count_29_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_29_load_0_req_1;
      LOAD_count_29_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_29_word_address_0;
      LOAD_count_29_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(69 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(319 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(94 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(4 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_start
  signal Block2_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_start
  signal Block3_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(18 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(10 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(0 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(4 downto 4),
      memory_space_3_sr_ack => memory_space_3_sr_ack(4 downto 4),
      memory_space_3_sr_addr => memory_space_3_sr_addr(69 downto 56),
      memory_space_3_sr_data => memory_space_3_sr_data(319 downto 256),
      memory_space_3_sr_tag => memory_space_3_sr_tag(94 downto 76),
      memory_space_3_sc_req => memory_space_3_sc_req(4 downto 4),
      memory_space_3_sc_ack => memory_space_3_sc_ack(4 downto 4),
      memory_space_3_sc_tag => memory_space_3_sc_tag(4 downto 4),
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(15 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(15 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(15 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(15 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(15 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(15 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(3 downto 3),
      memory_space_1_lr_ack => memory_space_1_lr_ack(3 downto 3),
      memory_space_1_lr_addr => memory_space_1_lr_addr(55 downto 42),
      memory_space_1_lr_tag => memory_space_1_lr_tag(75 downto 57),
      memory_space_1_lc_req => memory_space_1_lc_req(3 downto 3),
      memory_space_1_lc_ack => memory_space_1_lc_ack(3 downto 3),
      memory_space_1_lc_data => memory_space_1_lc_data(255 downto 192),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 3),
      memory_space_3_sr_req => memory_space_3_sr_req(3 downto 3),
      memory_space_3_sr_ack => memory_space_3_sr_ack(3 downto 3),
      memory_space_3_sr_addr => memory_space_3_sr_addr(55 downto 42),
      memory_space_3_sr_data => memory_space_3_sr_data(255 downto 192),
      memory_space_3_sr_tag => memory_space_3_sr_tag(75 downto 57),
      memory_space_3_sc_req => memory_space_3_sc_req(3 downto 3),
      memory_space_3_sc_ack => memory_space_3_sc_ack(3 downto 3),
      memory_space_3_sc_tag => memory_space_3_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(41 downto 28),
      memory_space_1_lr_tag => memory_space_1_lr_tag(56 downto 38),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(191 downto 128),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 2),
      memory_space_3_sr_req => memory_space_3_sr_req(2 downto 2),
      memory_space_3_sr_ack => memory_space_3_sr_ack(2 downto 2),
      memory_space_3_sr_addr => memory_space_3_sr_addr(41 downto 28),
      memory_space_3_sr_data => memory_space_3_sr_data(191 downto 128),
      memory_space_3_sr_tag => memory_space_3_sr_tag(56 downto 38),
      memory_space_3_sc_req => memory_space_3_sc_req(2 downto 2),
      memory_space_3_sc_ack => memory_space_3_sc_ack(2 downto 2),
      memory_space_3_sc_tag => memory_space_3_sc_tag(2 downto 2),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(15 downto 0),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(27 downto 14),
      memory_space_1_lr_tag => memory_space_1_lr_tag(37 downto 19),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(127 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 1),
      memory_space_3_sr_req => memory_space_3_sr_req(1 downto 1),
      memory_space_3_sr_ack => memory_space_3_sr_ack(1 downto 1),
      memory_space_3_sr_addr => memory_space_3_sr_addr(27 downto 14),
      memory_space_3_sr_data => memory_space_3_sr_data(127 downto 64),
      memory_space_3_sr_tag => memory_space_3_sr_tag(37 downto 19),
      memory_space_3_sc_req => memory_space_3_sc_req(1 downto 1),
      memory_space_3_sc_ack => memory_space_3_sc_ack(1 downto 1),
      memory_space_3_sc_tag => memory_space_3_sc_tag(1 downto 1),
      Block2_start_pipe_read_req => Block2_start_pipe_read_req(0 downto 0),
      Block2_start_pipe_read_ack => Block2_start_pipe_read_ack(0 downto 0),
      Block2_start_pipe_read_data => Block2_start_pipe_read_data(15 downto 0),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(13 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(63 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(18 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(0 downto 0),
      Block3_start_pipe_read_req => Block3_start_pipe_read_req(0 downto 0),
      Block3_start_pipe_read_ack => Block3_start_pipe_read_ack(0 downto 0),
      Block3_start_pipe_read_data => Block3_start_pipe_read_data(15 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(0 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(0 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  dummyROM_memory_space_0: dummy_read_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_2: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 1,
      num_stores => 5,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
