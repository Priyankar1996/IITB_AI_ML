-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_call_acks : in   std_logic_vector(0 downto 0);
    testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
    testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_return_acks : in   std_logic_vector(0 downto 0);
    testConfigure_return_data : in   std_logic_vector(15 downto 0);
    testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(31 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_call_acks : in   std_logic_vector(0 downto 0);
    sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
    sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_return_acks : in   std_logic_vector(0 downto 0);
    sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_4849_start: Boolean;
  signal convTranspose_CP_4849_symbol: Boolean;
  -- volatile/operator module components. 
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal WPIPE_Block1_start_1632_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_1645_inst_req_1 : boolean;
  signal call_stmt_1627_call_req_0 : boolean;
  signal call_stmt_1627_call_ack_0 : boolean;
  signal WPIPE_Block3_start_1640_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1632_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1632_inst_req_0 : boolean;
  signal call_stmt_1624_call_req_0 : boolean;
  signal call_stmt_1627_call_req_1 : boolean;
  signal call_stmt_1627_call_ack_1 : boolean;
  signal WPIPE_Block0_start_1628_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1632_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1640_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1640_inst_ack_0 : boolean;
  signal call_stmt_1624_call_ack_0 : boolean;
  signal RPIPE_Block1_done_1648_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1648_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_1645_inst_ack_1 : boolean;
  signal RPIPE_Block0_done_1645_inst_ack_0 : boolean;
  signal call_stmt_1624_call_req_1 : boolean;
  signal call_stmt_1624_call_ack_1 : boolean;
  signal RPIPE_Block0_done_1645_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1628_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1636_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1628_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1628_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1640_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1636_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1636_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1636_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1648_inst_req_1 : boolean;
  signal RPIPE_Block1_done_1648_inst_ack_1 : boolean;
  signal RPIPE_Block2_done_1651_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1651_inst_ack_0 : boolean;
  signal RPIPE_Block2_done_1651_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1651_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1654_inst_req_0 : boolean;
  signal RPIPE_Block3_done_1654_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1654_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1654_inst_ack_1 : boolean;
  signal call_stmt_1658_call_req_0 : boolean;
  signal call_stmt_1658_call_ack_0 : boolean;
  signal call_stmt_1658_call_req_1 : boolean;
  signal call_stmt_1658_call_ack_1 : boolean;
  signal type_cast_1666_inst_req_0 : boolean;
  signal type_cast_1666_inst_ack_0 : boolean;
  signal type_cast_1666_inst_req_1 : boolean;
  signal type_cast_1666_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1668_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1668_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1668_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1668_inst_ack_1 : boolean;
  signal call_stmt_1671_call_req_0 : boolean;
  signal call_stmt_1671_call_ack_0 : boolean;
  signal call_stmt_1671_call_req_1 : boolean;
  signal call_stmt_1671_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_4849_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_4849_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_4849_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_4849_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_4849: Block -- control-path 
    signal convTranspose_CP_4849_elements: BooleanArray(30 downto 0);
    -- 
  begin -- 
    convTranspose_CP_4849_elements(0) <= convTranspose_CP_4849_start;
    convTranspose_CP_4849_symbol <= convTranspose_CP_4849_elements(30);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 branch_block_stmt_1622/call_stmt_1624__entry__
      -- CP-element group 0: 	 branch_block_stmt_1622/call_stmt_1624/call_stmt_1624_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1622/call_stmt_1624/call_stmt_1624_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1622/call_stmt_1624/$entry
      -- CP-element group 0: 	 branch_block_stmt_1622/call_stmt_1624/call_stmt_1624_Sample/crr
      -- CP-element group 0: 	 branch_block_stmt_1622/call_stmt_1624/call_stmt_1624_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1622/call_stmt_1624/call_stmt_1624_Update/ccr
      -- CP-element group 0: 	 branch_block_stmt_1622/call_stmt_1624/call_stmt_1624_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1622/branch_block_stmt_1622__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1622/$entry
      -- 
    crr_4875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(0), ack => call_stmt_1624_call_req_0); -- 
    ccr_4880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(0), ack => call_stmt_1624_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_1622/call_stmt_1624/call_stmt_1624_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1622/call_stmt_1624/call_stmt_1624_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1622/call_stmt_1624/call_stmt_1624_Sample/cra
      -- 
    cra_4876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1624_call_ack_0, ack => convTranspose_CP_4849_elements(1)); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	9 
    -- CP-element group 2:  members (37) 
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1624__exit__
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655__entry__
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/call_stmt_1627_Sample/crr
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block0_done_1645_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block3_start_1640_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block1_start_1632_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1624/call_stmt_1624_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block1_done_1648_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block1_start_1632_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block3_start_1640_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/call_stmt_1627_Update/ccr
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block0_start_1628_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/call_stmt_1627_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block0_start_1628_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block1_start_1632_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block3_start_1640_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block1_done_1648_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block1_done_1648_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1624/call_stmt_1624_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1624/call_stmt_1624_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block2_start_1636_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1624/$exit
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block0_start_1628_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block0_done_1645_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/$entry
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/call_stmt_1627_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block0_done_1645_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/call_stmt_1627_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block2_start_1636_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block2_start_1636_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/call_stmt_1627_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block2_done_1651_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block2_done_1651_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block2_done_1651_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block3_done_1654_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block3_done_1654_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block3_done_1654_Sample/rr
      -- 
    cca_4881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1624_call_ack_1, ack => convTranspose_CP_4849_elements(2)); -- 
    crr_4892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(2), ack => call_stmt_1627_call_req_0); -- 
    req_4948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(2), ack => WPIPE_Block3_start_1640_inst_req_0); -- 
    req_4920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(2), ack => WPIPE_Block1_start_1632_inst_req_0); -- 
    ccr_4897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(2), ack => call_stmt_1627_call_req_1); -- 
    req_4906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(2), ack => WPIPE_Block0_start_1628_inst_req_0); -- 
    rr_4976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(2), ack => RPIPE_Block1_done_1648_inst_req_0); -- 
    rr_4962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(2), ack => RPIPE_Block0_done_1645_inst_req_0); -- 
    req_4934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(2), ack => WPIPE_Block2_start_1636_inst_req_0); -- 
    rr_4990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(2), ack => RPIPE_Block2_done_1651_inst_req_0); -- 
    rr_5004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(2), ack => RPIPE_Block3_done_1654_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/call_stmt_1627_Sample/cra
      -- CP-element group 3: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/call_stmt_1627_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/call_stmt_1627_sample_completed_
      -- 
    cra_4893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1627_call_ack_0, ack => convTranspose_CP_4849_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	21 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/call_stmt_1627_Update/cca
      -- CP-element group 4: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/call_stmt_1627_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/call_stmt_1627_update_completed_
      -- 
    cca_4898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1627_call_ack_1, ack => convTranspose_CP_4849_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block0_start_1628_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block0_start_1628_Sample/ack
      -- CP-element group 5: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block0_start_1628_Update/req
      -- CP-element group 5: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block0_start_1628_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block0_start_1628_update_start_
      -- CP-element group 5: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block0_start_1628_sample_completed_
      -- 
    ack_4907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1628_inst_ack_0, ack => convTranspose_CP_4849_elements(5)); -- 
    req_4911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(5), ack => WPIPE_Block0_start_1628_inst_req_1); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	21 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block0_start_1628_Update/ack
      -- CP-element group 6: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block0_start_1628_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block0_start_1628_update_completed_
      -- 
    ack_4912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1628_inst_ack_1, ack => convTranspose_CP_4849_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block1_start_1632_Sample/ack
      -- CP-element group 7: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block1_start_1632_Update/req
      -- CP-element group 7: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block1_start_1632_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block1_start_1632_update_start_
      -- CP-element group 7: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block1_start_1632_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block1_start_1632_Update/$entry
      -- 
    ack_4921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1632_inst_ack_0, ack => convTranspose_CP_4849_elements(7)); -- 
    req_4925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(7), ack => WPIPE_Block1_start_1632_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block1_start_1632_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block1_start_1632_Update/ack
      -- CP-element group 8: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block1_start_1632_update_completed_
      -- 
    ack_4926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1632_inst_ack_1, ack => convTranspose_CP_4849_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block2_start_1636_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block2_start_1636_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block2_start_1636_Update/req
      -- CP-element group 9: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block2_start_1636_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block2_start_1636_Sample/ack
      -- CP-element group 9: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block2_start_1636_Sample/$exit
      -- 
    ack_4935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1636_inst_ack_0, ack => convTranspose_CP_4849_elements(9)); -- 
    req_4939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(9), ack => WPIPE_Block2_start_1636_inst_req_1); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	21 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block2_start_1636_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block2_start_1636_Update/ack
      -- CP-element group 10: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block2_start_1636_Update/$exit
      -- 
    ack_4940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1636_inst_ack_1, ack => convTranspose_CP_4849_elements(10)); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block3_start_1640_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block3_start_1640_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block3_start_1640_update_start_
      -- CP-element group 11: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block3_start_1640_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block3_start_1640_Sample/ack
      -- CP-element group 11: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block3_start_1640_Update/req
      -- 
    ack_4949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1640_inst_ack_0, ack => convTranspose_CP_4849_elements(11)); -- 
    req_4953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(11), ack => WPIPE_Block3_start_1640_inst_req_1); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	21 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block3_start_1640_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block3_start_1640_Update/ack
      -- CP-element group 12: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/WPIPE_Block3_start_1640_Update/$exit
      -- 
    ack_4954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1640_inst_ack_1, ack => convTranspose_CP_4849_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block0_done_1645_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block0_done_1645_Update/cr
      -- CP-element group 13: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block0_done_1645_update_start_
      -- CP-element group 13: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block0_done_1645_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block0_done_1645_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block0_done_1645_Sample/ra
      -- 
    ra_4963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1645_inst_ack_0, ack => convTranspose_CP_4849_elements(13)); -- 
    cr_4967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(13), ack => RPIPE_Block0_done_1645_inst_req_1); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	21 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block0_done_1645_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block0_done_1645_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block0_done_1645_Update/ca
      -- 
    ca_4968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1645_inst_ack_1, ack => convTranspose_CP_4849_elements(14)); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block1_done_1648_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block1_done_1648_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block1_done_1648_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block1_done_1648_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block1_done_1648_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block1_done_1648_Update/cr
      -- 
    ra_4977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1648_inst_ack_0, ack => convTranspose_CP_4849_elements(15)); -- 
    cr_4981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(15), ack => RPIPE_Block1_done_1648_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	21 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block1_done_1648_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block1_done_1648_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block1_done_1648_Update/ca
      -- 
    ca_4982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1648_inst_ack_1, ack => convTranspose_CP_4849_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block2_done_1651_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block2_done_1651_update_start_
      -- CP-element group 17: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block2_done_1651_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block2_done_1651_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block2_done_1651_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block2_done_1651_Update/cr
      -- 
    ra_4991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1651_inst_ack_0, ack => convTranspose_CP_4849_elements(17)); -- 
    cr_4995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(17), ack => RPIPE_Block2_done_1651_inst_req_1); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block2_done_1651_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block2_done_1651_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block2_done_1651_Update/ca
      -- 
    ca_4996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1651_inst_ack_1, ack => convTranspose_CP_4849_elements(18)); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block3_done_1654_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block3_done_1654_update_start_
      -- CP-element group 19: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block3_done_1654_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block3_done_1654_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block3_done_1654_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block3_done_1654_Update/cr
      -- 
    ra_5005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1654_inst_ack_0, ack => convTranspose_CP_4849_elements(19)); -- 
    cr_5009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(19), ack => RPIPE_Block3_done_1654_inst_req_1); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block3_done_1654_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block3_done_1654_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/RPIPE_Block3_done_1654_Update/ca
      -- 
    ca_5010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1654_inst_ack_1, ack => convTranspose_CP_4849_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  place  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	12 
    -- CP-element group 21: 	16 
    -- CP-element group 21: 	18 
    -- CP-element group 21: 	20 
    -- CP-element group 21: 	6 
    -- CP-element group 21: 	4 
    -- CP-element group 21: 	14 
    -- CP-element group 21: 	8 
    -- CP-element group 21: 	10 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	23 
    -- CP-element group 21: 	25 
    -- CP-element group 21: 	28 
    -- CP-element group 21: 	29 
    -- CP-element group 21:  members (19) 
      -- CP-element group 21: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671__entry__
      -- CP-element group 21: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655__exit__
      -- CP-element group 21: 	 branch_block_stmt_1622/call_stmt_1627_to_assign_stmt_1655/$exit
      -- CP-element group 21: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/$entry
      -- CP-element group 21: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1658_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1658_update_start_
      -- CP-element group 21: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1658_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1658_Sample/crr
      -- CP-element group 21: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1658_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1658_Update/ccr
      -- CP-element group 21: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/type_cast_1666_update_start_
      -- CP-element group 21: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/type_cast_1666_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/type_cast_1666_Update/cr
      -- CP-element group 21: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1671_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1671_update_start_
      -- CP-element group 21: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1671_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1671_Sample/crr
      -- CP-element group 21: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1671_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1671_Update/ccr
      -- 
    crr_5021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(21), ack => call_stmt_1658_call_req_0); -- 
    ccr_5026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(21), ack => call_stmt_1658_call_req_1); -- 
    cr_5040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(21), ack => type_cast_1666_inst_req_1); -- 
    crr_5063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(21), ack => call_stmt_1671_call_req_0); -- 
    ccr_5068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(21), ack => call_stmt_1671_call_req_1); -- 
    convTranspose_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_4849_elements(12) & convTranspose_CP_4849_elements(16) & convTranspose_CP_4849_elements(18) & convTranspose_CP_4849_elements(20) & convTranspose_CP_4849_elements(6) & convTranspose_CP_4849_elements(4) & convTranspose_CP_4849_elements(14) & convTranspose_CP_4849_elements(8) & convTranspose_CP_4849_elements(10);
      gj_convTranspose_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_4849_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1658_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1658_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1658_Sample/cra
      -- 
    cra_5022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1658_call_ack_0, ack => convTranspose_CP_4849_elements(22)); -- 
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1658_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1658_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1658_Update/cca
      -- CP-element group 23: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/type_cast_1666_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/type_cast_1666_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/type_cast_1666_Sample/rr
      -- 
    cca_5027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1658_call_ack_1, ack => convTranspose_CP_4849_elements(23)); -- 
    rr_5035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(23), ack => type_cast_1666_inst_req_0); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/type_cast_1666_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/type_cast_1666_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/type_cast_1666_Sample/ra
      -- 
    ra_5036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1666_inst_ack_0, ack => convTranspose_CP_4849_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	21 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/type_cast_1666_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/type_cast_1666_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/type_cast_1666_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/WPIPE_elapsed_time_pipe_1668_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/WPIPE_elapsed_time_pipe_1668_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/WPIPE_elapsed_time_pipe_1668_Sample/req
      -- 
    ca_5041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1666_inst_ack_1, ack => convTranspose_CP_4849_elements(25)); -- 
    req_5049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(25), ack => WPIPE_elapsed_time_pipe_1668_inst_req_0); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/WPIPE_elapsed_time_pipe_1668_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/WPIPE_elapsed_time_pipe_1668_update_start_
      -- CP-element group 26: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/WPIPE_elapsed_time_pipe_1668_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/WPIPE_elapsed_time_pipe_1668_Sample/ack
      -- CP-element group 26: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/WPIPE_elapsed_time_pipe_1668_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/WPIPE_elapsed_time_pipe_1668_Update/req
      -- 
    ack_5050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1668_inst_ack_0, ack => convTranspose_CP_4849_elements(26)); -- 
    req_5054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_4849_elements(26), ack => WPIPE_elapsed_time_pipe_1668_inst_req_1); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	30 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/WPIPE_elapsed_time_pipe_1668_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/WPIPE_elapsed_time_pipe_1668_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/WPIPE_elapsed_time_pipe_1668_Update/ack
      -- 
    ack_5055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1668_inst_ack_1, ack => convTranspose_CP_4849_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	21 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1671_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1671_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1671_Sample/cra
      -- 
    cra_5064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1671_call_ack_0, ack => convTranspose_CP_4849_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	21 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1671_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1671_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/call_stmt_1671_Update/cca
      -- 
    cca_5069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1671_call_ack_1, ack => convTranspose_CP_4849_elements(29)); -- 
    -- CP-element group 30:  join  transition  place  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (13) 
      -- CP-element group 30: 	 branch_block_stmt_1622/branch_block_stmt_1622__exit__
      -- CP-element group 30: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671__exit__
      -- CP-element group 30: 	 branch_block_stmt_1622/return__
      -- CP-element group 30: 	 branch_block_stmt_1622/merge_stmt_1673__exit__
      -- CP-element group 30: 	 $exit
      -- CP-element group 30: 	 branch_block_stmt_1622/$exit
      -- CP-element group 30: 	 branch_block_stmt_1622/call_stmt_1658_to_call_stmt_1671/$exit
      -- CP-element group 30: 	 branch_block_stmt_1622/return___PhiReq/$entry
      -- CP-element group 30: 	 branch_block_stmt_1622/return___PhiReq/$exit
      -- CP-element group 30: 	 branch_block_stmt_1622/merge_stmt_1673_PhiReqMerge
      -- CP-element group 30: 	 branch_block_stmt_1622/merge_stmt_1673_PhiAck/$entry
      -- CP-element group 30: 	 branch_block_stmt_1622/merge_stmt_1673_PhiAck/$exit
      -- CP-element group 30: 	 branch_block_stmt_1622/merge_stmt_1673_PhiAck/dummy
      -- 
    convTranspose_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_4849_elements(27) & convTranspose_CP_4849_elements(29);
      gj_convTranspose_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_4849_elements(30), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal call10_1652 : std_logic_vector(15 downto 0);
    signal call12_1655 : std_logic_vector(15 downto 0);
    signal call14_1658 : std_logic_vector(31 downto 0);
    signal call1_1627 : std_logic_vector(31 downto 0);
    signal call6_1646 : std_logic_vector(15 downto 0);
    signal call8_1649 : std_logic_vector(15 downto 0);
    signal call_1624 : std_logic_vector(15 downto 0);
    signal conv_1667 : std_logic_vector(63 downto 0);
    signal sub_1663 : std_logic_vector(31 downto 0);
    signal type_cast_1630_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1634_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1638_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1642_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    type_cast_1630_wire_constant <= "0000000000000001";
    type_cast_1634_wire_constant <= "0000000000000001";
    type_cast_1638_wire_constant <= "0000000000000001";
    type_cast_1642_wire_constant <= "0000000000000001";
    type_cast_1666_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1666_inst_req_0;
      type_cast_1666_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1666_inst_req_1;
      type_cast_1666_inst_ack_1<= rack(0);
      type_cast_1666_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1666_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_1663,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1667,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- binary operator SUB_u32_u32_1662_inst
    process(call14_1658, call1_1627) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(call14_1658, call1_1627, tmp_var);
      sub_1663 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_Block0_done_1645_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1645_inst_req_0;
      RPIPE_Block0_done_1645_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1645_inst_req_1;
      RPIPE_Block0_done_1645_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call6_1646 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1648_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1648_inst_req_0;
      RPIPE_Block1_done_1648_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1648_inst_req_1;
      RPIPE_Block1_done_1648_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call8_1649 <= data_out(15 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1651_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1651_inst_req_0;
      RPIPE_Block2_done_1651_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1651_inst_req_1;
      RPIPE_Block2_done_1651_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call10_1652 <= data_out(15 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1654_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1654_inst_req_0;
      RPIPE_Block3_done_1654_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1654_inst_req_1;
      RPIPE_Block3_done_1654_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call12_1655 <= data_out(15 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_Block0_start_1628_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_start_1628_inst_req_0;
      WPIPE_Block0_start_1628_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_start_1628_inst_req_1;
      WPIPE_Block0_start_1628_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1630_wire_constant;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_1632_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_start_1632_inst_req_0;
      WPIPE_Block1_start_1632_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_start_1632_inst_req_1;
      WPIPE_Block1_start_1632_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1634_wire_constant;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1636_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_start_1636_inst_req_0;
      WPIPE_Block2_start_1636_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_start_1636_inst_req_1;
      WPIPE_Block2_start_1636_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1638_wire_constant;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1640_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_start_1640_inst_req_0;
      WPIPE_Block3_start_1640_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_start_1640_inst_req_1;
      WPIPE_Block3_start_1640_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1642_wire_constant;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_elapsed_time_pipe_1668_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1668_inst_req_0;
      WPIPE_elapsed_time_pipe_1668_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1668_inst_req_1;
      WPIPE_elapsed_time_pipe_1668_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= conv_1667;
      elapsed_time_pipe_write_4_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_4: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared call operator group (0) : call_stmt_1624_call 
    testConfigure_call_group_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1624_call_req_0;
      call_stmt_1624_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1624_call_req_1;
      call_stmt_1624_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      testConfigure_call_group_0_gI: SplitGuardInterface generic map(name => "testConfigure_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call_1624 <= data_out(15 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => testConfigure_call_reqs(0),
          ackR => testConfigure_call_acks(0),
          tagR => testConfigure_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 16,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => testConfigure_return_acks(0), -- cross-over
          ackL => testConfigure_return_reqs(0), -- cross-over
          dataL => testConfigure_return_data(15 downto 0),
          tagL => testConfigure_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1627_call call_stmt_1658_call 
    timer_call_group_1: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1627_call_req_0;
      reqL_unguarded(0) <= call_stmt_1658_call_req_0;
      call_stmt_1627_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1658_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1627_call_req_1;
      reqR_unguarded(0) <= call_stmt_1658_call_req_1;
      call_stmt_1627_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1658_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_1_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_1_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_1_gI: SplitGuardInterface generic map(name => "timer_call_group_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call1_1627 <= data_out(63 downto 32);
      call14_1658 <= data_out(31 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(31 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1671_call 
    sendOutput_call_group_2: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1671_call_req_0;
      call_stmt_1671_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1671_call_req_1;
      call_stmt_1671_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendOutput_call_group_2_gI: SplitGuardInterface generic map(name => "sendOutput_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => sendOutput_call_reqs(0),
          ackR => sendOutput_call_acks(0),
          tagR => sendOutput_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendOutput_return_acks(0), -- cross-over
          ackL => sendOutput_return_reqs(0), -- cross-over
          tagL => sendOutput_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_5078_start: Boolean;
  signal convTransposeA_CP_5078_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1946_inst_req_1 : boolean;
  signal addr_of_1983_final_reg_ack_1 : boolean;
  signal addr_of_1953_final_reg_req_1 : boolean;
  signal type_cast_1946_inst_ack_1 : boolean;
  signal addr_of_1953_final_reg_ack_1 : boolean;
  signal array_obj_ref_1982_index_offset_req_0 : boolean;
  signal addr_of_1983_final_reg_req_1 : boolean;
  signal type_cast_1962_inst_req_0 : boolean;
  signal type_cast_1976_inst_ack_0 : boolean;
  signal array_obj_ref_1982_index_offset_ack_0 : boolean;
  signal type_cast_1962_inst_ack_0 : boolean;
  signal array_obj_ref_1982_index_offset_req_1 : boolean;
  signal type_cast_1976_inst_req_1 : boolean;
  signal ptr_deref_1801_load_0_req_1 : boolean;
  signal ptr_deref_1801_load_0_ack_1 : boolean;
  signal type_cast_1976_inst_req_0 : boolean;
  signal array_obj_ref_1982_index_offset_ack_1 : boolean;
  signal ptr_deref_1957_load_0_req_1 : boolean;
  signal addr_of_1983_final_reg_req_0 : boolean;
  signal addr_of_1983_final_reg_ack_0 : boolean;
  signal type_cast_1976_inst_ack_1 : boolean;
  signal type_cast_1805_inst_req_0 : boolean;
  signal type_cast_1962_inst_req_1 : boolean;
  signal type_cast_1962_inst_ack_1 : boolean;
  signal ptr_deref_1957_load_0_req_0 : boolean;
  signal ptr_deref_1957_load_0_ack_0 : boolean;
  signal ptr_deref_1986_store_0_req_0 : boolean;
  signal ptr_deref_1986_store_0_ack_0 : boolean;
  signal array_obj_ref_1952_index_offset_req_0 : boolean;
  signal array_obj_ref_1952_index_offset_ack_0 : boolean;
  signal ptr_deref_1957_load_0_ack_1 : boolean;
  signal RPIPE_Block0_start_1679_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1679_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1679_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1679_inst_ack_1 : boolean;
  signal type_cast_1946_inst_ack_0 : boolean;
  signal type_cast_1946_inst_req_0 : boolean;
  signal addr_of_1953_final_reg_ack_0 : boolean;
  signal addr_of_1953_final_reg_req_0 : boolean;
  signal ptr_deref_1801_load_0_ack_0 : boolean;
  signal ptr_deref_1692_load_0_req_0 : boolean;
  signal ptr_deref_1692_load_0_ack_0 : boolean;
  signal ptr_deref_1692_load_0_req_1 : boolean;
  signal type_cast_1931_inst_ack_1 : boolean;
  signal ptr_deref_1692_load_0_ack_1 : boolean;
  signal type_cast_1931_inst_req_1 : boolean;
  signal ptr_deref_1801_load_0_req_0 : boolean;
  signal type_cast_1931_inst_ack_0 : boolean;
  signal type_cast_1931_inst_req_0 : boolean;
  signal ptr_deref_1704_load_0_req_0 : boolean;
  signal ptr_deref_1704_load_0_ack_0 : boolean;
  signal ptr_deref_1704_load_0_req_1 : boolean;
  signal ptr_deref_1704_load_0_ack_1 : boolean;
  signal array_obj_ref_1952_index_offset_ack_1 : boolean;
  signal type_cast_1805_inst_ack_1 : boolean;
  signal type_cast_1805_inst_req_1 : boolean;
  signal array_obj_ref_1952_index_offset_req_1 : boolean;
  signal type_cast_1805_inst_ack_0 : boolean;
  signal ptr_deref_1714_load_0_req_0 : boolean;
  signal ptr_deref_1714_load_0_ack_0 : boolean;
  signal ptr_deref_1714_load_0_req_1 : boolean;
  signal ptr_deref_1714_load_0_ack_1 : boolean;
  signal ptr_deref_1726_load_0_req_0 : boolean;
  signal ptr_deref_1726_load_0_ack_0 : boolean;
  signal ptr_deref_1726_load_0_req_1 : boolean;
  signal ptr_deref_1726_load_0_ack_1 : boolean;
  signal LOAD_padding_1729_load_0_req_0 : boolean;
  signal LOAD_padding_1729_load_0_ack_0 : boolean;
  signal LOAD_padding_1729_load_0_req_1 : boolean;
  signal LOAD_padding_1729_load_0_ack_1 : boolean;
  signal ptr_deref_1739_load_0_req_0 : boolean;
  signal ptr_deref_1739_load_0_ack_0 : boolean;
  signal ptr_deref_1739_load_0_req_1 : boolean;
  signal ptr_deref_1739_load_0_ack_1 : boolean;
  signal ptr_deref_1751_load_0_req_0 : boolean;
  signal ptr_deref_1751_load_0_ack_0 : boolean;
  signal ptr_deref_1751_load_0_req_1 : boolean;
  signal ptr_deref_1751_load_0_ack_1 : boolean;
  signal ptr_deref_1763_load_0_req_0 : boolean;
  signal ptr_deref_1763_load_0_ack_0 : boolean;
  signal ptr_deref_1763_load_0_req_1 : boolean;
  signal ptr_deref_1763_load_0_ack_1 : boolean;
  signal ptr_deref_1775_load_0_req_0 : boolean;
  signal ptr_deref_1775_load_0_ack_0 : boolean;
  signal ptr_deref_1775_load_0_req_1 : boolean;
  signal ptr_deref_1775_load_0_ack_1 : boolean;
  signal type_cast_1779_inst_req_0 : boolean;
  signal type_cast_1779_inst_ack_0 : boolean;
  signal type_cast_1779_inst_req_1 : boolean;
  signal type_cast_1779_inst_ack_1 : boolean;
  signal type_cast_1783_inst_req_0 : boolean;
  signal type_cast_1783_inst_ack_0 : boolean;
  signal type_cast_1783_inst_req_1 : boolean;
  signal type_cast_1783_inst_ack_1 : boolean;
  signal ptr_deref_1986_store_0_req_1 : boolean;
  signal ptr_deref_1986_store_0_ack_1 : boolean;
  signal type_cast_1992_inst_req_0 : boolean;
  signal type_cast_1992_inst_ack_0 : boolean;
  signal type_cast_1992_inst_req_1 : boolean;
  signal type_cast_1992_inst_ack_1 : boolean;
  signal if_stmt_2007_branch_req_0 : boolean;
  signal if_stmt_2007_branch_ack_1 : boolean;
  signal if_stmt_2007_branch_ack_0 : boolean;
  signal type_cast_2031_inst_req_0 : boolean;
  signal type_cast_2031_inst_ack_0 : boolean;
  signal type_cast_2031_inst_req_1 : boolean;
  signal type_cast_2031_inst_ack_1 : boolean;
  signal type_cast_2040_inst_req_0 : boolean;
  signal type_cast_2040_inst_ack_0 : boolean;
  signal type_cast_2040_inst_req_1 : boolean;
  signal type_cast_2040_inst_ack_1 : boolean;
  signal type_cast_2057_inst_req_0 : boolean;
  signal type_cast_2057_inst_ack_0 : boolean;
  signal type_cast_2057_inst_req_1 : boolean;
  signal type_cast_2057_inst_ack_1 : boolean;
  signal if_stmt_2064_branch_req_0 : boolean;
  signal if_stmt_2064_branch_ack_1 : boolean;
  signal if_stmt_2064_branch_ack_0 : boolean;
  signal WPIPE_Block0_done_2072_inst_req_0 : boolean;
  signal WPIPE_Block0_done_2072_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_2072_inst_req_1 : boolean;
  signal WPIPE_Block0_done_2072_inst_ack_1 : boolean;
  signal phi_stmt_1844_req_0 : boolean;
  signal phi_stmt_1837_req_0 : boolean;
  signal type_cast_1850_inst_req_0 : boolean;
  signal type_cast_1850_inst_ack_0 : boolean;
  signal type_cast_1850_inst_req_1 : boolean;
  signal type_cast_1850_inst_ack_1 : boolean;
  signal phi_stmt_1844_req_1 : boolean;
  signal type_cast_1843_inst_req_0 : boolean;
  signal type_cast_1843_inst_ack_0 : boolean;
  signal type_cast_1843_inst_req_1 : boolean;
  signal type_cast_1843_inst_ack_1 : boolean;
  signal phi_stmt_1837_req_1 : boolean;
  signal phi_stmt_1837_ack_0 : boolean;
  signal phi_stmt_1844_ack_0 : boolean;
  signal type_cast_1907_inst_req_0 : boolean;
  signal type_cast_1907_inst_ack_0 : boolean;
  signal type_cast_1907_inst_req_1 : boolean;
  signal type_cast_1907_inst_ack_1 : boolean;
  signal phi_stmt_1904_req_0 : boolean;
  signal phi_stmt_1904_req_1 : boolean;
  signal phi_stmt_1904_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_5078_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_5078_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_5078_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_5078_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_5078: Block -- control-path 
    signal convTransposeA_CP_5078_elements: BooleanArray(85 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_5078_elements(0) <= convTransposeA_CP_5078_start;
    convTransposeA_CP_5078_symbol <= convTransposeA_CP_5078_elements(65);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1677/$entry
      -- CP-element group 0: 	 branch_block_stmt_1677/branch_block_stmt_1677__entry__
      -- CP-element group 0: 	 branch_block_stmt_1677/assign_stmt_1680__entry__
      -- CP-element group 0: 	 branch_block_stmt_1677/assign_stmt_1680/$entry
      -- CP-element group 0: 	 branch_block_stmt_1677/assign_stmt_1680/RPIPE_Block0_start_1679_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1677/assign_stmt_1680/RPIPE_Block0_start_1679_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1677/assign_stmt_1680/RPIPE_Block0_start_1679_Sample/rr
      -- 
    rr_5126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(0), ack => RPIPE_Block0_start_1679_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1677/assign_stmt_1680/RPIPE_Block0_start_1679_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1677/assign_stmt_1680/RPIPE_Block0_start_1679_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1677/assign_stmt_1680/RPIPE_Block0_start_1679_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1677/assign_stmt_1680/RPIPE_Block0_start_1679_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1677/assign_stmt_1680/RPIPE_Block0_start_1679_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1677/assign_stmt_1680/RPIPE_Block0_start_1679_Update/cr
      -- 
    ra_5127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1679_inst_ack_0, ack => convTransposeA_CP_5078_elements(1)); -- 
    cr_5131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(1), ack => RPIPE_Block0_start_1679_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	25 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (262) 
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1680__exit__
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834__entry__
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1680/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1680/RPIPE_Block0_start_1679_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1680/RPIPE_Block0_start_1679_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1680/RPIPE_Block0_start_1679_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1805_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1805_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1805_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1779_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1779_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1779_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1783_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1783_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1783_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_base_address_calculated
      -- 
    ca_5132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1679_inst_ack_1, ack => convTransposeA_CP_5078_elements(2)); -- 
    cr_5640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => ptr_deref_1801_load_0_req_1); -- 
    rr_5168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => ptr_deref_1692_load_0_req_0); -- 
    cr_5179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => ptr_deref_1692_load_0_req_1); -- 
    rr_5629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => ptr_deref_1801_load_0_req_0); -- 
    rr_5218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => ptr_deref_1704_load_0_req_0); -- 
    cr_5229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => ptr_deref_1704_load_0_req_1); -- 
    cr_5659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => type_cast_1805_inst_req_1); -- 
    rr_5268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => ptr_deref_1714_load_0_req_0); -- 
    cr_5279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => ptr_deref_1714_load_0_req_1); -- 
    rr_5318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => ptr_deref_1726_load_0_req_0); -- 
    cr_5329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => ptr_deref_1726_load_0_req_1); -- 
    rr_5351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => LOAD_padding_1729_load_0_req_0); -- 
    cr_5362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => LOAD_padding_1729_load_0_req_1); -- 
    rr_5401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => ptr_deref_1739_load_0_req_0); -- 
    cr_5412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => ptr_deref_1739_load_0_req_1); -- 
    rr_5451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => ptr_deref_1751_load_0_req_0); -- 
    cr_5462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => ptr_deref_1751_load_0_req_1); -- 
    rr_5501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => ptr_deref_1763_load_0_req_0); -- 
    cr_5512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => ptr_deref_1763_load_0_req_1); -- 
    rr_5551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => ptr_deref_1775_load_0_req_0); -- 
    cr_5562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => ptr_deref_1775_load_0_req_1); -- 
    cr_5581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => type_cast_1779_inst_req_1); -- 
    cr_5595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(2), ack => type_cast_1783_inst_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_Sample/word_access_start/word_0/ra
      -- 
    ra_5169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1692_load_0_ack_0, ack => convTransposeA_CP_5078_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	21 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_Update/ptr_deref_1692_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_Update/ptr_deref_1692_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_Update/ptr_deref_1692_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1692_Update/ptr_deref_1692_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1779_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1779_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1779_Sample/rr
      -- 
    ca_5180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1692_load_0_ack_1, ack => convTransposeA_CP_5078_elements(4)); -- 
    rr_5576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(4), ack => type_cast_1779_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_Sample/word_access_start/word_0/ra
      -- 
    ra_5219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1704_load_0_ack_0, ack => convTransposeA_CP_5078_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	23 
    -- CP-element group 6:  members (12) 
      -- CP-element group 6: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_Update/ptr_deref_1704_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_Update/ptr_deref_1704_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_Update/ptr_deref_1704_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1704_Update/ptr_deref_1704_Merge/merge_ack
      -- CP-element group 6: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1783_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1783_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1783_Sample/rr
      -- 
    ca_5230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1704_load_0_ack_1, ack => convTransposeA_CP_5078_elements(6)); -- 
    rr_5590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(6), ack => type_cast_1783_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_Sample/word_access_start/word_0/ra
      -- 
    ra_5269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1714_load_0_ack_0, ack => convTransposeA_CP_5078_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	29 
    -- CP-element group 8:  members (9) 
      -- CP-element group 8: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_Update/ptr_deref_1714_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_Update/ptr_deref_1714_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_Update/ptr_deref_1714_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1714_Update/ptr_deref_1714_Merge/merge_ack
      -- 
    ca_5280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1714_load_0_ack_1, ack => convTransposeA_CP_5078_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_Sample/word_access_start/word_0/ra
      -- 
    ra_5319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1726_load_0_ack_0, ack => convTransposeA_CP_5078_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	29 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_Update/ptr_deref_1726_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_Update/ptr_deref_1726_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_Update/ptr_deref_1726_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1726_Update/ptr_deref_1726_Merge/merge_ack
      -- 
    ca_5330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1726_load_0_ack_1, ack => convTransposeA_CP_5078_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_Sample/word_access_start/word_0/ra
      -- 
    ra_5352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1729_load_0_ack_0, ack => convTransposeA_CP_5078_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	29 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_Update/LOAD_padding_1729_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_Update/LOAD_padding_1729_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_Update/LOAD_padding_1729_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/LOAD_padding_1729_Update/LOAD_padding_1729_Merge/merge_ack
      -- 
    ca_5363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1729_load_0_ack_1, ack => convTransposeA_CP_5078_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_Sample/word_access_start/word_0/ra
      -- 
    ra_5402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1739_load_0_ack_0, ack => convTransposeA_CP_5078_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	29 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_Update/ptr_deref_1739_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_Update/ptr_deref_1739_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_Update/ptr_deref_1739_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1739_Update/ptr_deref_1739_Merge/merge_ack
      -- 
    ca_5413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1739_load_0_ack_1, ack => convTransposeA_CP_5078_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_Sample/word_access_start/word_0/ra
      -- 
    ra_5452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1751_load_0_ack_0, ack => convTransposeA_CP_5078_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	29 
    -- CP-element group 16:  members (9) 
      -- CP-element group 16: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_Update/ptr_deref_1751_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_Update/ptr_deref_1751_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_Update/ptr_deref_1751_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1751_Update/ptr_deref_1751_Merge/merge_ack
      -- 
    ca_5463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1751_load_0_ack_1, ack => convTransposeA_CP_5078_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_Sample/word_access_start/word_0/ra
      -- 
    ra_5502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1763_load_0_ack_0, ack => convTransposeA_CP_5078_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	29 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_Update/ptr_deref_1763_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_Update/ptr_deref_1763_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_Update/ptr_deref_1763_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1763_Update/ptr_deref_1763_Merge/merge_ack
      -- 
    ca_5513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1763_load_0_ack_1, ack => convTransposeA_CP_5078_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_Sample/word_access_start/word_0/ra
      -- 
    ra_5552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1775_load_0_ack_0, ack => convTransposeA_CP_5078_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	29 
    -- CP-element group 20:  members (9) 
      -- CP-element group 20: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_Update/ptr_deref_1775_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_Update/ptr_deref_1775_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_Update/ptr_deref_1775_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1775_Update/ptr_deref_1775_Merge/merge_ack
      -- 
    ca_5563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1775_load_0_ack_1, ack => convTransposeA_CP_5078_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	4 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1779_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1779_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1779_Sample/ra
      -- 
    ra_5577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1779_inst_ack_0, ack => convTransposeA_CP_5078_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	29 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1779_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1779_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1779_Update/ca
      -- 
    ca_5582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1779_inst_ack_1, ack => convTransposeA_CP_5078_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	6 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1783_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1783_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1783_Sample/ra
      -- 
    ra_5591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1783_inst_ack_0, ack => convTransposeA_CP_5078_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	29 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1783_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1783_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1783_Update/ca
      -- 
    ca_5596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1783_inst_ack_1, ack => convTransposeA_CP_5078_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_Sample/word_access_start/word_0/ra
      -- CP-element group 25: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_sample_completed_
      -- 
    ra_5630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1801_load_0_ack_0, ack => convTransposeA_CP_5078_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (12) 
      -- CP-element group 26: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_Update/word_access_complete/word_0/ca
      -- CP-element group 26: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_Update/ptr_deref_1801_Merge/$entry
      -- CP-element group 26: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_Update/ptr_deref_1801_Merge/$exit
      -- CP-element group 26: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_Update/ptr_deref_1801_Merge/merge_req
      -- CP-element group 26: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1805_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1805_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1805_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_Update/ptr_deref_1801_Merge/merge_ack
      -- CP-element group 26: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/ptr_deref_1801_update_completed_
      -- 
    ca_5641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1801_load_0_ack_1, ack => convTransposeA_CP_5078_elements(26)); -- 
    rr_5654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(26), ack => type_cast_1805_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1805_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1805_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1805_Sample/ra
      -- 
    ra_5655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1805_inst_ack_0, ack => convTransposeA_CP_5078_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1805_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1805_Update/ca
      -- CP-element group 28: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/type_cast_1805_Update/$exit
      -- 
    ca_5660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1805_inst_ack_1, ack => convTransposeA_CP_5078_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  place  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	8 
    -- CP-element group 29: 	16 
    -- CP-element group 29: 	18 
    -- CP-element group 29: 	20 
    -- CP-element group 29: 	22 
    -- CP-element group 29: 	24 
    -- CP-element group 29: 	28 
    -- CP-element group 29: 	10 
    -- CP-element group 29: 	12 
    -- CP-element group 29: 	14 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	66 
    -- CP-element group 29: 	67 
    -- CP-element group 29:  members (8) 
      -- CP-element group 29: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834__exit__
      -- CP-element group 29: 	 branch_block_stmt_1677/entry_whilex_xbodyx_xouter
      -- CP-element group 29: 	 branch_block_stmt_1677/assign_stmt_1689_to_assign_stmt_1834/$exit
      -- CP-element group 29: 	 branch_block_stmt_1677/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 29: 	 branch_block_stmt_1677/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/$entry
      -- CP-element group 29: 	 branch_block_stmt_1677/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/phi_stmt_1844_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_1677/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/$entry
      -- CP-element group 29: 	 branch_block_stmt_1677/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/phi_stmt_1837_sources/$entry
      -- 
    convTransposeA_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeA_CP_5078_elements(8) & convTransposeA_CP_5078_elements(16) & convTransposeA_CP_5078_elements(18) & convTransposeA_CP_5078_elements(20) & convTransposeA_CP_5078_elements(22) & convTransposeA_CP_5078_elements(24) & convTransposeA_CP_5078_elements(28) & convTransposeA_CP_5078_elements(10) & convTransposeA_CP_5078_elements(12) & convTransposeA_CP_5078_elements(14);
      gj_convTransposeA_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_5078_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	85 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1931_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1931_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1931_sample_completed_
      -- 
    ra_5675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1931_inst_ack_0, ack => convTransposeA_CP_5078_elements(30)); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	85 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1946_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1946_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1946_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1931_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1931_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1931_update_completed_
      -- 
    ca_5680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1931_inst_ack_1, ack => convTransposeA_CP_5078_elements(31)); -- 
    rr_5688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(31), ack => type_cast_1946_inst_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1946_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1946_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1946_sample_completed_
      -- 
    ra_5689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1946_inst_ack_0, ack => convTransposeA_CP_5078_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	85 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (16) 
      -- CP-element group 33: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1946_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_index_resized_1
      -- CP-element group 33: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_index_scaled_1
      -- CP-element group 33: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_index_computed_1
      -- CP-element group 33: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_index_resize_1/$entry
      -- CP-element group 33: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_final_index_sum_regn_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_index_resize_1/$exit
      -- CP-element group 33: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_index_resize_1/index_resize_req
      -- CP-element group 33: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_final_index_sum_regn_Sample/req
      -- CP-element group 33: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_index_resize_1/index_resize_ack
      -- CP-element group 33: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_index_scale_1/$entry
      -- CP-element group 33: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_index_scale_1/$exit
      -- CP-element group 33: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_index_scale_1/scale_rename_req
      -- CP-element group 33: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_index_scale_1/scale_rename_ack
      -- CP-element group 33: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1946_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1946_update_completed_
      -- 
    ca_5694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1946_inst_ack_1, ack => convTransposeA_CP_5078_elements(33)); -- 
    req_5719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(33), ack => array_obj_ref_1952_index_offset_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	53 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_final_index_sum_regn_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_final_index_sum_regn_Sample/ack
      -- CP-element group 34: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_final_index_sum_regn_sample_complete
      -- 
    ack_5720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1952_index_offset_ack_0, ack => convTransposeA_CP_5078_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	85 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (11) 
      -- CP-element group 35: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1953_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_root_address_calculated
      -- CP-element group 35: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_offset_calculated
      -- CP-element group 35: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_final_index_sum_regn_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1953_request/req
      -- CP-element group 35: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1953_request/$entry
      -- CP-element group 35: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_base_plus_offset/sum_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_base_plus_offset/sum_rename_req
      -- CP-element group 35: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_base_plus_offset/$exit
      -- CP-element group 35: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_base_plus_offset/$entry
      -- CP-element group 35: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_final_index_sum_regn_Update/ack
      -- 
    ack_5725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1952_index_offset_ack_1, ack => convTransposeA_CP_5078_elements(35)); -- 
    req_5734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(35), ack => addr_of_1953_final_reg_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1953_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1953_request/ack
      -- CP-element group 36: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1953_request/$exit
      -- 
    ack_5735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1953_final_reg_ack_0, ack => convTransposeA_CP_5078_elements(36)); -- 
    -- CP-element group 37:  join  fork  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	85 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (24) 
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1953_complete/$exit
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1953_complete/ack
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_word_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_word_addrgen/$entry
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_word_addrgen/$exit
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_word_addrgen/root_register_req
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_word_addrgen/root_register_ack
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_Sample/word_access_start/word_0/$entry
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_base_addr_resize/base_resize_req
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_base_addr_resize/base_resize_ack
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_base_plus_offset/$entry
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_Sample/word_access_start/word_0/rr
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1953_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_base_address_resized
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_base_addr_resize/$entry
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_base_addr_resize/$exit
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_base_plus_offset/sum_rename_req
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_base_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_base_plus_offset/$exit
      -- CP-element group 37: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_Sample/word_access_start/$entry
      -- 
    ack_5740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1953_final_reg_ack_1, ack => convTransposeA_CP_5078_elements(37)); -- 
    rr_5773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(37), ack => ptr_deref_1957_load_0_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_Sample/word_access_start/word_0/$exit
      -- CP-element group 38: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_Sample/word_access_start/word_0/ra
      -- CP-element group 38: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_Sample/word_access_start/$exit
      -- 
    ra_5774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1957_load_0_ack_0, ack => convTransposeA_CP_5078_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	85 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	48 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_Update/word_access_complete/word_0/$exit
      -- CP-element group 39: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_Update/ptr_deref_1957_Merge/$entry
      -- CP-element group 39: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_Update/ptr_deref_1957_Merge/merge_req
      -- CP-element group 39: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_Update/ptr_deref_1957_Merge/$exit
      -- CP-element group 39: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_Update/ptr_deref_1957_Merge/merge_ack
      -- CP-element group 39: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_Update/word_access_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_Update/word_access_complete/word_0/ca
      -- CP-element group 39: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_update_completed_
      -- 
    ca_5785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1957_load_0_ack_1, ack => convTransposeA_CP_5078_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	85 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1962_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1962_Sample/ra
      -- CP-element group 40: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1962_sample_completed_
      -- 
    ra_5799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1962_inst_ack_0, ack => convTransposeA_CP_5078_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	85 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1962_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1976_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1976_Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1962_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1962_Update/ca
      -- CP-element group 41: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1976_sample_start_
      -- 
    ca_5804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1962_inst_ack_1, ack => convTransposeA_CP_5078_elements(41)); -- 
    rr_5812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(41), ack => type_cast_1976_inst_req_0); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1976_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1976_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1976_sample_completed_
      -- 
    ra_5813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1976_inst_ack_0, ack => convTransposeA_CP_5078_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	85 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (16) 
      -- CP-element group 43: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_final_index_sum_regn_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_final_index_sum_regn_Sample/req
      -- CP-element group 43: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1976_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1976_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1976_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_index_resize_1/$entry
      -- CP-element group 43: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_index_resize_1/$exit
      -- CP-element group 43: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_index_resize_1/index_resize_req
      -- CP-element group 43: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_index_resize_1/index_resize_ack
      -- CP-element group 43: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_index_resized_1
      -- CP-element group 43: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_index_scaled_1
      -- CP-element group 43: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_index_scale_1/$exit
      -- CP-element group 43: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_index_computed_1
      -- CP-element group 43: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_index_scale_1/scale_rename_req
      -- CP-element group 43: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_index_scale_1/scale_rename_ack
      -- CP-element group 43: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_index_scale_1/$entry
      -- 
    ca_5818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1976_inst_ack_1, ack => convTransposeA_CP_5078_elements(43)); -- 
    req_5843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(43), ack => array_obj_ref_1982_index_offset_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	53 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_final_index_sum_regn_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_final_index_sum_regn_sample_complete
      -- CP-element group 44: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_final_index_sum_regn_Sample/ack
      -- 
    ack_5844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1982_index_offset_ack_0, ack => convTransposeA_CP_5078_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	85 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (11) 
      -- CP-element group 45: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_final_index_sum_regn_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_final_index_sum_regn_Update/ack
      -- CP-element group 45: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_base_plus_offset/$entry
      -- CP-element group 45: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_base_plus_offset/$exit
      -- CP-element group 45: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_base_plus_offset/sum_rename_req
      -- CP-element group 45: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_base_plus_offset/sum_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1983_request/$entry
      -- CP-element group 45: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1983_request/req
      -- CP-element group 45: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_root_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1983_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_offset_calculated
      -- 
    ack_5849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1982_index_offset_ack_1, ack => convTransposeA_CP_5078_elements(45)); -- 
    req_5858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(45), ack => addr_of_1983_final_reg_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1983_request/$exit
      -- CP-element group 46: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1983_request/ack
      -- CP-element group 46: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1983_sample_completed_
      -- 
    ack_5859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1983_final_reg_ack_0, ack => convTransposeA_CP_5078_elements(46)); -- 
    -- CP-element group 47:  fork  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	85 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (19) 
      -- CP-element group 47: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1983_complete/ack
      -- CP-element group 47: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_base_plus_offset/sum_rename_req
      -- CP-element group 47: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_word_addrgen/root_register_req
      -- CP-element group 47: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_base_plus_offset/sum_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_word_addrgen/$entry
      -- CP-element group 47: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_word_addrgen/$exit
      -- CP-element group 47: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1983_complete/$exit
      -- CP-element group 47: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_base_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1983_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_root_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_word_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_word_addrgen/root_register_ack
      -- CP-element group 47: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_base_plus_offset/$exit
      -- CP-element group 47: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_base_address_resized
      -- CP-element group 47: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_base_addr_resize/$entry
      -- CP-element group 47: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_base_addr_resize/$exit
      -- CP-element group 47: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_base_addr_resize/base_resize_req
      -- CP-element group 47: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_base_addr_resize/base_resize_ack
      -- CP-element group 47: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_base_plus_offset/$entry
      -- 
    ack_5864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1983_final_reg_ack_1, ack => convTransposeA_CP_5078_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	39 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (9) 
      -- CP-element group 48: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_Sample/ptr_deref_1986_Split/$entry
      -- CP-element group 48: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_Sample/ptr_deref_1986_Split/$exit
      -- CP-element group 48: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_Sample/ptr_deref_1986_Split/split_req
      -- CP-element group 48: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_Sample/ptr_deref_1986_Split/split_ack
      -- CP-element group 48: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_Sample/word_access_start/word_0/rr
      -- CP-element group 48: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_Sample/word_access_start/word_0/$entry
      -- CP-element group 48: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_Sample/word_access_start/$entry
      -- 
    rr_5902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(48), ack => ptr_deref_1986_store_0_req_0); -- 
    convTransposeA_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_5078_elements(39) & convTransposeA_CP_5078_elements(47);
      gj_convTransposeA_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_5078_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_Sample/word_access_start/$exit
      -- CP-element group 49: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_Sample/word_access_start/word_0/ra
      -- CP-element group 49: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_Sample/word_access_start/word_0/$exit
      -- 
    ra_5903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1986_store_0_ack_0, ack => convTransposeA_CP_5078_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	85 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_Update/word_access_complete/word_0/$exit
      -- CP-element group 50: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_Update/word_access_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_Update/word_access_complete/word_0/ca
      -- 
    ca_5914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1986_store_0_ack_1, ack => convTransposeA_CP_5078_elements(50)); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	85 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1992_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1992_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1992_Sample/ra
      -- 
    ra_5923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1992_inst_ack_0, ack => convTransposeA_CP_5078_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	85 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1992_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1992_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1992_Update/ca
      -- 
    ca_5928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1992_inst_ack_1, ack => convTransposeA_CP_5078_elements(52)); -- 
    -- CP-element group 53:  branch  join  transition  place  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	34 
    -- CP-element group 53: 	44 
    -- CP-element group 53: 	50 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (10) 
      -- CP-element group 53: 	 branch_block_stmt_1677/R_cmp_2008_place
      -- CP-element group 53: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006__exit__
      -- CP-element group 53: 	 branch_block_stmt_1677/if_stmt_2007__entry__
      -- CP-element group 53: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/$exit
      -- CP-element group 53: 	 branch_block_stmt_1677/if_stmt_2007_dead_link/$entry
      -- CP-element group 53: 	 branch_block_stmt_1677/if_stmt_2007_eval_test/$entry
      -- CP-element group 53: 	 branch_block_stmt_1677/if_stmt_2007_eval_test/$exit
      -- CP-element group 53: 	 branch_block_stmt_1677/if_stmt_2007_eval_test/branch_req
      -- CP-element group 53: 	 branch_block_stmt_1677/if_stmt_2007_if_link/$entry
      -- CP-element group 53: 	 branch_block_stmt_1677/if_stmt_2007_else_link/$entry
      -- 
    branch_req_5936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(53), ack => if_stmt_2007_branch_req_0); -- 
    convTransposeA_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_5078_elements(34) & convTransposeA_CP_5078_elements(44) & convTransposeA_CP_5078_elements(50) & convTransposeA_CP_5078_elements(52);
      gj_convTransposeA_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_5078_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	80 
    -- CP-element group 54: 	81 
    -- CP-element group 54:  members (24) 
      -- CP-element group 54: 	 branch_block_stmt_1677/whilex_xbody_ifx_xthen
      -- CP-element group 54: 	 branch_block_stmt_1677/merge_stmt_2013__exit__
      -- CP-element group 54: 	 branch_block_stmt_1677/assign_stmt_2019__entry__
      -- CP-element group 54: 	 branch_block_stmt_1677/assign_stmt_2019__exit__
      -- CP-element group 54: 	 branch_block_stmt_1677/ifx_xthen_whilex_xbody
      -- CP-element group 54: 	 branch_block_stmt_1677/if_stmt_2007_if_link/$exit
      -- CP-element group 54: 	 branch_block_stmt_1677/if_stmt_2007_if_link/if_choice_transition
      -- CP-element group 54: 	 branch_block_stmt_1677/assign_stmt_2019/$entry
      -- CP-element group 54: 	 branch_block_stmt_1677/assign_stmt_2019/$exit
      -- CP-element group 54: 	 branch_block_stmt_1677/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_1677/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1904/$entry
      -- CP-element group 54: 	 branch_block_stmt_1677/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1904/phi_stmt_1904_sources/$entry
      -- CP-element group 54: 	 branch_block_stmt_1677/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1904/phi_stmt_1904_sources/type_cast_1907/$entry
      -- CP-element group 54: 	 branch_block_stmt_1677/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1904/phi_stmt_1904_sources/type_cast_1907/SplitProtocol/$entry
      -- CP-element group 54: 	 branch_block_stmt_1677/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1904/phi_stmt_1904_sources/type_cast_1907/SplitProtocol/Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_1677/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1904/phi_stmt_1904_sources/type_cast_1907/SplitProtocol/Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_1677/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1904/phi_stmt_1904_sources/type_cast_1907/SplitProtocol/Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_1677/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1904/phi_stmt_1904_sources/type_cast_1907/SplitProtocol/Update/cr
      -- CP-element group 54: 	 branch_block_stmt_1677/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_1677/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 54: 	 branch_block_stmt_1677/merge_stmt_2013_PhiReqMerge
      -- CP-element group 54: 	 branch_block_stmt_1677/merge_stmt_2013_PhiAck/$entry
      -- CP-element group 54: 	 branch_block_stmt_1677/merge_stmt_2013_PhiAck/$exit
      -- CP-element group 54: 	 branch_block_stmt_1677/merge_stmt_2013_PhiAck/dummy
      -- 
    if_choice_transition_5941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2007_branch_ack_1, ack => convTransposeA_CP_5078_elements(54)); -- 
    rr_6124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(54), ack => type_cast_1907_inst_req_0); -- 
    cr_6129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(54), ack => type_cast_1907_inst_req_1); -- 
    -- CP-element group 55:  fork  transition  place  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	57 
    -- CP-element group 55: 	59 
    -- CP-element group 55: 	61 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_1677/whilex_xbody_ifx_xelse
      -- CP-element group 55: 	 branch_block_stmt_1677/merge_stmt_2021__exit__
      -- CP-element group 55: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063__entry__
      -- CP-element group 55: 	 branch_block_stmt_1677/if_stmt_2007_else_link/$exit
      -- CP-element group 55: 	 branch_block_stmt_1677/if_stmt_2007_else_link/else_choice_transition
      -- CP-element group 55: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/$entry
      -- CP-element group 55: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2031_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2031_update_start_
      -- CP-element group 55: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2031_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2031_Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2031_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2031_Update/cr
      -- CP-element group 55: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2040_update_start_
      -- CP-element group 55: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2040_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2040_Update/cr
      -- CP-element group 55: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2057_update_start_
      -- CP-element group 55: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2057_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2057_Update/cr
      -- CP-element group 55: 	 branch_block_stmt_1677/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 55: 	 branch_block_stmt_1677/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 55: 	 branch_block_stmt_1677/merge_stmt_2021_PhiReqMerge
      -- CP-element group 55: 	 branch_block_stmt_1677/merge_stmt_2021_PhiAck/$entry
      -- CP-element group 55: 	 branch_block_stmt_1677/merge_stmt_2021_PhiAck/$exit
      -- CP-element group 55: 	 branch_block_stmt_1677/merge_stmt_2021_PhiAck/dummy
      -- 
    else_choice_transition_5945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2007_branch_ack_0, ack => convTransposeA_CP_5078_elements(55)); -- 
    rr_5961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(55), ack => type_cast_2031_inst_req_0); -- 
    cr_5966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(55), ack => type_cast_2031_inst_req_1); -- 
    cr_5980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(55), ack => type_cast_2040_inst_req_1); -- 
    cr_5994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(55), ack => type_cast_2057_inst_req_1); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2031_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2031_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2031_Sample/ra
      -- 
    ra_5962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2031_inst_ack_0, ack => convTransposeA_CP_5078_elements(56)); -- 
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2031_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2031_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2031_Update/ca
      -- CP-element group 57: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2040_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2040_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2040_Sample/rr
      -- 
    ca_5967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2031_inst_ack_1, ack => convTransposeA_CP_5078_elements(57)); -- 
    rr_5975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(57), ack => type_cast_2040_inst_req_0); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2040_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2040_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2040_Sample/ra
      -- 
    ra_5976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2040_inst_ack_0, ack => convTransposeA_CP_5078_elements(58)); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	55 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2040_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2040_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2040_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2057_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2057_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2057_Sample/rr
      -- 
    ca_5981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2040_inst_ack_1, ack => convTransposeA_CP_5078_elements(59)); -- 
    rr_5989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(59), ack => type_cast_2057_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2057_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2057_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2057_Sample/ra
      -- 
    ra_5990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2057_inst_ack_0, ack => convTransposeA_CP_5078_elements(60)); -- 
    -- CP-element group 61:  branch  transition  place  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	55 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (13) 
      -- CP-element group 61: 	 branch_block_stmt_1677/R_cmp86_2065_place
      -- CP-element group 61: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063__exit__
      -- CP-element group 61: 	 branch_block_stmt_1677/if_stmt_2064__entry__
      -- CP-element group 61: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/$exit
      -- CP-element group 61: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2057_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2057_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_1677/assign_stmt_2027_to_assign_stmt_2063/type_cast_2057_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_1677/if_stmt_2064_dead_link/$entry
      -- CP-element group 61: 	 branch_block_stmt_1677/if_stmt_2064_eval_test/$entry
      -- CP-element group 61: 	 branch_block_stmt_1677/if_stmt_2064_eval_test/$exit
      -- CP-element group 61: 	 branch_block_stmt_1677/if_stmt_2064_eval_test/branch_req
      -- CP-element group 61: 	 branch_block_stmt_1677/if_stmt_2064_if_link/$entry
      -- CP-element group 61: 	 branch_block_stmt_1677/if_stmt_2064_else_link/$entry
      -- 
    ca_5995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2057_inst_ack_1, ack => convTransposeA_CP_5078_elements(61)); -- 
    branch_req_6003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(61), ack => if_stmt_2064_branch_req_0); -- 
    -- CP-element group 62:  merge  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (15) 
      -- CP-element group 62: 	 branch_block_stmt_1677/ifx_xelse_whilex_xend
      -- CP-element group 62: 	 branch_block_stmt_1677/merge_stmt_2070__exit__
      -- CP-element group 62: 	 branch_block_stmt_1677/assign_stmt_2074__entry__
      -- CP-element group 62: 	 branch_block_stmt_1677/if_stmt_2064_if_link/$exit
      -- CP-element group 62: 	 branch_block_stmt_1677/if_stmt_2064_if_link/if_choice_transition
      -- CP-element group 62: 	 branch_block_stmt_1677/assign_stmt_2074/$entry
      -- CP-element group 62: 	 branch_block_stmt_1677/assign_stmt_2074/WPIPE_Block0_done_2072_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1677/assign_stmt_2074/WPIPE_Block0_done_2072_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1677/assign_stmt_2074/WPIPE_Block0_done_2072_Sample/req
      -- CP-element group 62: 	 branch_block_stmt_1677/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 62: 	 branch_block_stmt_1677/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 62: 	 branch_block_stmt_1677/merge_stmt_2070_PhiReqMerge
      -- CP-element group 62: 	 branch_block_stmt_1677/merge_stmt_2070_PhiAck/$entry
      -- CP-element group 62: 	 branch_block_stmt_1677/merge_stmt_2070_PhiAck/$exit
      -- CP-element group 62: 	 branch_block_stmt_1677/merge_stmt_2070_PhiAck/dummy
      -- 
    if_choice_transition_6008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2064_branch_ack_1, ack => convTransposeA_CP_5078_elements(62)); -- 
    req_6025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(62), ack => WPIPE_Block0_done_2072_inst_req_0); -- 
    -- CP-element group 63:  fork  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	69 
    -- CP-element group 63: 	70 
    -- CP-element group 63: 	72 
    -- CP-element group 63: 	73 
    -- CP-element group 63:  members (20) 
      -- CP-element group 63: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 63: 	 branch_block_stmt_1677/if_stmt_2064_else_link/$exit
      -- CP-element group 63: 	 branch_block_stmt_1677/if_stmt_2064_else_link/else_choice_transition
      -- CP-element group 63: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 63: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/$entry
      -- CP-element group 63: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/phi_stmt_1844_sources/$entry
      -- CP-element group 63: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/phi_stmt_1844_sources/type_cast_1850/$entry
      -- CP-element group 63: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/phi_stmt_1844_sources/type_cast_1850/SplitProtocol/$entry
      -- CP-element group 63: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/phi_stmt_1844_sources/type_cast_1850/SplitProtocol/Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/phi_stmt_1844_sources/type_cast_1850/SplitProtocol/Sample/rr
      -- CP-element group 63: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/phi_stmt_1844_sources/type_cast_1850/SplitProtocol/Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/phi_stmt_1844_sources/type_cast_1850/SplitProtocol/Update/cr
      -- CP-element group 63: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/$entry
      -- CP-element group 63: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/phi_stmt_1837_sources/$entry
      -- CP-element group 63: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/phi_stmt_1837_sources/type_cast_1843/$entry
      -- CP-element group 63: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/phi_stmt_1837_sources/type_cast_1843/SplitProtocol/$entry
      -- CP-element group 63: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/phi_stmt_1837_sources/type_cast_1843/SplitProtocol/Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/phi_stmt_1837_sources/type_cast_1843/SplitProtocol/Sample/rr
      -- CP-element group 63: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/phi_stmt_1837_sources/type_cast_1843/SplitProtocol/Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/phi_stmt_1837_sources/type_cast_1843/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2064_branch_ack_0, ack => convTransposeA_CP_5078_elements(63)); -- 
    rr_6069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(63), ack => type_cast_1850_inst_req_0); -- 
    cr_6074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(63), ack => type_cast_1850_inst_req_1); -- 
    rr_6092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(63), ack => type_cast_1843_inst_req_0); -- 
    cr_6097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(63), ack => type_cast_1843_inst_req_1); -- 
    -- CP-element group 64:  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (6) 
      -- CP-element group 64: 	 branch_block_stmt_1677/assign_stmt_2074/WPIPE_Block0_done_2072_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1677/assign_stmt_2074/WPIPE_Block0_done_2072_update_start_
      -- CP-element group 64: 	 branch_block_stmt_1677/assign_stmt_2074/WPIPE_Block0_done_2072_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1677/assign_stmt_2074/WPIPE_Block0_done_2072_Sample/ack
      -- CP-element group 64: 	 branch_block_stmt_1677/assign_stmt_2074/WPIPE_Block0_done_2072_Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_1677/assign_stmt_2074/WPIPE_Block0_done_2072_Update/req
      -- 
    ack_6026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_2072_inst_ack_0, ack => convTransposeA_CP_5078_elements(64)); -- 
    req_6030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(64), ack => WPIPE_Block0_done_2072_inst_req_1); -- 
    -- CP-element group 65:  transition  place  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (16) 
      -- CP-element group 65: 	 $exit
      -- CP-element group 65: 	 branch_block_stmt_1677/$exit
      -- CP-element group 65: 	 branch_block_stmt_1677/branch_block_stmt_1677__exit__
      -- CP-element group 65: 	 branch_block_stmt_1677/assign_stmt_2074__exit__
      -- CP-element group 65: 	 branch_block_stmt_1677/return__
      -- CP-element group 65: 	 branch_block_stmt_1677/merge_stmt_2076__exit__
      -- CP-element group 65: 	 branch_block_stmt_1677/assign_stmt_2074/$exit
      -- CP-element group 65: 	 branch_block_stmt_1677/assign_stmt_2074/WPIPE_Block0_done_2072_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1677/assign_stmt_2074/WPIPE_Block0_done_2072_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1677/assign_stmt_2074/WPIPE_Block0_done_2072_Update/ack
      -- CP-element group 65: 	 branch_block_stmt_1677/return___PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_1677/return___PhiReq/$exit
      -- CP-element group 65: 	 branch_block_stmt_1677/merge_stmt_2076_PhiReqMerge
      -- CP-element group 65: 	 branch_block_stmt_1677/merge_stmt_2076_PhiAck/$entry
      -- CP-element group 65: 	 branch_block_stmt_1677/merge_stmt_2076_PhiAck/$exit
      -- CP-element group 65: 	 branch_block_stmt_1677/merge_stmt_2076_PhiAck/dummy
      -- 
    ack_6031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_2072_inst_ack_1, ack => convTransposeA_CP_5078_elements(65)); -- 
    -- CP-element group 66:  transition  output  delay-element  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	29 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_1677/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/$exit
      -- CP-element group 66: 	 branch_block_stmt_1677/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/phi_stmt_1844_sources/$exit
      -- CP-element group 66: 	 branch_block_stmt_1677/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/phi_stmt_1844_sources/type_cast_1848_konst_delay_trans
      -- CP-element group 66: 	 branch_block_stmt_1677/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/phi_stmt_1844_req
      -- 
    phi_stmt_1844_req_6042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1844_req_6042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(66), ack => phi_stmt_1844_req_0); -- 
    -- Element group convTransposeA_CP_5078_elements(66) is a control-delay.
    cp_element_66_delay: control_delay_element  generic map(name => " 66_delay", delay_value => 1)  port map(req => convTransposeA_CP_5078_elements(29), ack => convTransposeA_CP_5078_elements(66), clk => clk, reset =>reset);
    -- CP-element group 67:  transition  output  delay-element  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	29 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_1677/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/$exit
      -- CP-element group 67: 	 branch_block_stmt_1677/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/phi_stmt_1837_sources/$exit
      -- CP-element group 67: 	 branch_block_stmt_1677/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/phi_stmt_1837_sources/type_cast_1841_konst_delay_trans
      -- CP-element group 67: 	 branch_block_stmt_1677/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/phi_stmt_1837_req
      -- 
    phi_stmt_1837_req_6050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1837_req_6050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(67), ack => phi_stmt_1837_req_0); -- 
    -- Element group convTransposeA_CP_5078_elements(67) is a control-delay.
    cp_element_67_delay: control_delay_element  generic map(name => " 67_delay", delay_value => 1)  port map(req => convTransposeA_CP_5078_elements(29), ack => convTransposeA_CP_5078_elements(67), clk => clk, reset =>reset);
    -- CP-element group 68:  join  transition  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	76 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_1677/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_5078_elements(66) & convTransposeA_CP_5078_elements(67);
      gj_convTransposeA_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_5078_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	63 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/phi_stmt_1844_sources/type_cast_1850/SplitProtocol/Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/phi_stmt_1844_sources/type_cast_1850/SplitProtocol/Sample/ra
      -- 
    ra_6070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1850_inst_ack_0, ack => convTransposeA_CP_5078_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	63 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/phi_stmt_1844_sources/type_cast_1850/SplitProtocol/Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/phi_stmt_1844_sources/type_cast_1850/SplitProtocol/Update/ca
      -- 
    ca_6075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1850_inst_ack_1, ack => convTransposeA_CP_5078_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	75 
    -- CP-element group 71:  members (5) 
      -- CP-element group 71: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/$exit
      -- CP-element group 71: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/phi_stmt_1844_sources/$exit
      -- CP-element group 71: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/phi_stmt_1844_sources/type_cast_1850/$exit
      -- CP-element group 71: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/phi_stmt_1844_sources/type_cast_1850/SplitProtocol/$exit
      -- CP-element group 71: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1844/phi_stmt_1844_req
      -- 
    phi_stmt_1844_req_6076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1844_req_6076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(71), ack => phi_stmt_1844_req_1); -- 
    convTransposeA_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_5078_elements(69) & convTransposeA_CP_5078_elements(70);
      gj_convTransposeA_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_5078_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	63 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/phi_stmt_1837_sources/type_cast_1843/SplitProtocol/Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/phi_stmt_1837_sources/type_cast_1843/SplitProtocol/Sample/ra
      -- 
    ra_6093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1843_inst_ack_0, ack => convTransposeA_CP_5078_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	63 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/phi_stmt_1837_sources/type_cast_1843/SplitProtocol/Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/phi_stmt_1837_sources/type_cast_1843/SplitProtocol/Update/ca
      -- 
    ca_6098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1843_inst_ack_1, ack => convTransposeA_CP_5078_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/$exit
      -- CP-element group 74: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/phi_stmt_1837_sources/$exit
      -- CP-element group 74: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/phi_stmt_1837_sources/type_cast_1843/$exit
      -- CP-element group 74: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/phi_stmt_1837_sources/type_cast_1843/SplitProtocol/$exit
      -- CP-element group 74: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1837/phi_stmt_1837_req
      -- 
    phi_stmt_1837_req_6099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1837_req_6099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(74), ack => phi_stmt_1837_req_1); -- 
    convTransposeA_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_5078_elements(72) & convTransposeA_CP_5078_elements(73);
      gj_convTransposeA_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_5078_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	71 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_1677/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_5078_elements(71) & convTransposeA_CP_5078_elements(74);
      gj_convTransposeA_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_5078_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  merge  fork  transition  place  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	68 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_1677/merge_stmt_1836_PhiReqMerge
      -- CP-element group 76: 	 branch_block_stmt_1677/merge_stmt_1836_PhiAck/$entry
      -- 
    convTransposeA_CP_5078_elements(76) <= OrReduce(convTransposeA_CP_5078_elements(68) & convTransposeA_CP_5078_elements(75));
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1677/merge_stmt_1836_PhiAck/phi_stmt_1837_ack
      -- 
    phi_stmt_1837_ack_6104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1837_ack_0, ack => convTransposeA_CP_5078_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1677/merge_stmt_1836_PhiAck/phi_stmt_1844_ack
      -- 
    phi_stmt_1844_ack_6105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1844_ack_0, ack => convTransposeA_CP_5078_elements(78)); -- 
    -- CP-element group 79:  join  transition  place  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	83 
    -- CP-element group 79:  members (10) 
      -- CP-element group 79: 	 branch_block_stmt_1677/merge_stmt_1836__exit__
      -- CP-element group 79: 	 branch_block_stmt_1677/assign_stmt_1856_to_assign_stmt_1901__entry__
      -- CP-element group 79: 	 branch_block_stmt_1677/assign_stmt_1856_to_assign_stmt_1901__exit__
      -- CP-element group 79: 	 branch_block_stmt_1677/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 79: 	 branch_block_stmt_1677/assign_stmt_1856_to_assign_stmt_1901/$exit
      -- CP-element group 79: 	 branch_block_stmt_1677/assign_stmt_1856_to_assign_stmt_1901/$entry
      -- CP-element group 79: 	 branch_block_stmt_1677/merge_stmt_1836_PhiAck/$exit
      -- CP-element group 79: 	 branch_block_stmt_1677/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 79: 	 branch_block_stmt_1677/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1904/$entry
      -- CP-element group 79: 	 branch_block_stmt_1677/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1904/phi_stmt_1904_sources/$entry
      -- 
    convTransposeA_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_5078_elements(77) & convTransposeA_CP_5078_elements(78);
      gj_convTransposeA_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_5078_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	54 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1677/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1904/phi_stmt_1904_sources/type_cast_1907/SplitProtocol/Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_1677/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1904/phi_stmt_1904_sources/type_cast_1907/SplitProtocol/Sample/ra
      -- 
    ra_6125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1907_inst_ack_0, ack => convTransposeA_CP_5078_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	54 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1677/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1904/phi_stmt_1904_sources/type_cast_1907/SplitProtocol/Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_1677/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1904/phi_stmt_1904_sources/type_cast_1907/SplitProtocol/Update/ca
      -- 
    ca_6130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1907_inst_ack_1, ack => convTransposeA_CP_5078_elements(81)); -- 
    -- CP-element group 82:  join  transition  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_1677/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 82: 	 branch_block_stmt_1677/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1904/$exit
      -- CP-element group 82: 	 branch_block_stmt_1677/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1904/phi_stmt_1904_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_1677/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1904/phi_stmt_1904_sources/type_cast_1907/$exit
      -- CP-element group 82: 	 branch_block_stmt_1677/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1904/phi_stmt_1904_sources/type_cast_1907/SplitProtocol/$exit
      -- CP-element group 82: 	 branch_block_stmt_1677/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1904/phi_stmt_1904_req
      -- 
    phi_stmt_1904_req_6131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1904_req_6131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(82), ack => phi_stmt_1904_req_0); -- 
    convTransposeA_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_5078_elements(80) & convTransposeA_CP_5078_elements(81);
      gj_convTransposeA_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_5078_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  transition  output  delay-element  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	79 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (5) 
      -- CP-element group 83: 	 branch_block_stmt_1677/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 83: 	 branch_block_stmt_1677/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1904/$exit
      -- CP-element group 83: 	 branch_block_stmt_1677/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1904/phi_stmt_1904_sources/$exit
      -- CP-element group 83: 	 branch_block_stmt_1677/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1904/phi_stmt_1904_sources/type_cast_1910_konst_delay_trans
      -- CP-element group 83: 	 branch_block_stmt_1677/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1904/phi_stmt_1904_req
      -- 
    phi_stmt_1904_req_6142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1904_req_6142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(83), ack => phi_stmt_1904_req_1); -- 
    -- Element group convTransposeA_CP_5078_elements(83) is a control-delay.
    cp_element_83_delay: control_delay_element  generic map(name => " 83_delay", delay_value => 1)  port map(req => convTransposeA_CP_5078_elements(79), ack => convTransposeA_CP_5078_elements(83), clk => clk, reset =>reset);
    -- CP-element group 84:  merge  transition  place  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1677/merge_stmt_1903_PhiReqMerge
      -- CP-element group 84: 	 branch_block_stmt_1677/merge_stmt_1903_PhiAck/$entry
      -- 
    convTransposeA_CP_5078_elements(84) <= OrReduce(convTransposeA_CP_5078_elements(82) & convTransposeA_CP_5078_elements(83));
    -- CP-element group 85:  fork  transition  place  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	30 
    -- CP-element group 85: 	31 
    -- CP-element group 85: 	33 
    -- CP-element group 85: 	35 
    -- CP-element group 85: 	37 
    -- CP-element group 85: 	39 
    -- CP-element group 85: 	40 
    -- CP-element group 85: 	41 
    -- CP-element group 85: 	43 
    -- CP-element group 85: 	45 
    -- CP-element group 85: 	47 
    -- CP-element group 85: 	50 
    -- CP-element group 85: 	51 
    -- CP-element group 85: 	52 
    -- CP-element group 85:  members (51) 
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1946_Update/cr
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1953_complete/req
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1962_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_final_index_sum_regn_update_start
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1983_complete/req
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1962_Sample/rr
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1983_complete/$entry
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_final_index_sum_regn_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_final_index_sum_regn_Update/req
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1976_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1976_Update/cr
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_Update/word_access_complete/word_0/cr
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1962_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1982_final_index_sum_regn_update_start
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_Update/word_access_complete/word_0/$entry
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1962_Update/cr
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1953_update_start_
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_update_start_
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_update_start_
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1962_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_Update/word_access_complete/$entry
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1983_update_start_
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1962_update_start_
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1976_update_start_
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_final_index_sum_regn_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_Update/word_access_complete/$entry
      -- CP-element group 85: 	 branch_block_stmt_1677/merge_stmt_1903__exit__
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006__entry__
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1957_Update/word_access_complete/word_0/$entry
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/addr_of_1953_complete/$entry
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1946_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1946_update_start_
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1931_Update/cr
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1931_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1931_Sample/rr
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1931_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1931_update_start_
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1931_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/$entry
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/array_obj_ref_1952_final_index_sum_regn_Update/req
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/ptr_deref_1986_Update/word_access_complete/word_0/cr
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1992_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1992_update_start_
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1992_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1992_Sample/rr
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1992_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_1677/assign_stmt_1917_to_assign_stmt_2006/type_cast_1992_Update/cr
      -- CP-element group 85: 	 branch_block_stmt_1677/merge_stmt_1903_PhiAck/$exit
      -- CP-element group 85: 	 branch_block_stmt_1677/merge_stmt_1903_PhiAck/phi_stmt_1904_ack
      -- 
    phi_stmt_1904_ack_6147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1904_ack_0, ack => convTransposeA_CP_5078_elements(85)); -- 
    cr_5693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(85), ack => type_cast_1946_inst_req_1); -- 
    req_5739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(85), ack => addr_of_1953_final_reg_req_1); -- 
    req_5863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(85), ack => addr_of_1983_final_reg_req_1); -- 
    rr_5798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(85), ack => type_cast_1962_inst_req_0); -- 
    req_5848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(85), ack => array_obj_ref_1982_index_offset_req_1); -- 
    cr_5817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(85), ack => type_cast_1976_inst_req_1); -- 
    cr_5784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(85), ack => ptr_deref_1957_load_0_req_1); -- 
    cr_5803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(85), ack => type_cast_1962_inst_req_1); -- 
    cr_5679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(85), ack => type_cast_1931_inst_req_1); -- 
    rr_5674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(85), ack => type_cast_1931_inst_req_0); -- 
    req_5724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(85), ack => array_obj_ref_1952_index_offset_req_1); -- 
    cr_5913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(85), ack => ptr_deref_1986_store_0_req_1); -- 
    rr_5922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(85), ack => type_cast_1992_inst_req_0); -- 
    cr_5927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_5078_elements(85), ack => type_cast_1992_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1939_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1970_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_1729_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_1729_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom58_1981_resized : std_logic_vector(13 downto 0);
    signal R_idxprom58_1981_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1951_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1951_scaled : std_logic_vector(13 downto 0);
    signal add10_1922 : std_logic_vector(15 downto 0);
    signal add50_1927 : std_logic_vector(15 downto 0);
    signal add63_1999 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1952_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1952_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1952_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1952_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1952_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1952_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1982_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1982_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1982_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1982_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1982_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1982_root_address : std_logic_vector(13 downto 0);
    signal arrayidx59_1984 : std_logic_vector(31 downto 0);
    signal arrayidx_1954 : std_logic_vector(31 downto 0);
    signal call_1680 : std_logic_vector(15 downto 0);
    signal cmp76_2037 : std_logic_vector(0 downto 0);
    signal cmp86_2063 : std_logic_vector(0 downto 0);
    signal cmp_2006 : std_logic_vector(0 downto 0);
    signal conv53_1932 : std_logic_vector(31 downto 0);
    signal conv56_1963 : std_logic_vector(31 downto 0);
    signal conv62_1993 : std_logic_vector(31 downto 0);
    signal conv65_1780 : std_logic_vector(31 downto 0);
    signal conv73_2032 : std_logic_vector(31 downto 0);
    signal conv75_1784 : std_logic_vector(31 downto 0);
    signal conv82_2058 : std_logic_vector(31 downto 0);
    signal conv84_1806 : std_logic_vector(31 downto 0);
    signal div85_1812 : std_logic_vector(31 downto 0);
    signal div_1790 : std_logic_vector(31 downto 0);
    signal iNsTr_10_1798 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1689 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1701 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1711 : std_logic_vector(31 downto 0);
    signal iNsTr_5_1723 : std_logic_vector(31 downto 0);
    signal iNsTr_6_1736 : std_logic_vector(31 downto 0);
    signal iNsTr_7_1748 : std_logic_vector(31 downto 0);
    signal iNsTr_8_1760 : std_logic_vector(31 downto 0);
    signal iNsTr_9_1772 : std_logic_vector(31 downto 0);
    signal idxprom58_1977 : std_logic_vector(63 downto 0);
    signal idxprom_1947 : std_logic_vector(63 downto 0);
    signal inc80_2041 : std_logic_vector(15 downto 0);
    signal inc80x_xinput_dim0x_x2_2046 : std_logic_vector(15 downto 0);
    signal inc_2027 : std_logic_vector(15 downto 0);
    signal indvar_1904 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2019 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_1844 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_1837 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2053 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1917 : std_logic_vector(15 downto 0);
    signal ptr_deref_1692_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1692_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1692_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1692_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1692_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1704_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1704_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1704_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1704_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1704_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1714_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1714_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1714_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1714_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1714_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1726_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1726_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1726_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1726_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1726_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1739_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1739_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1739_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1739_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1739_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1751_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1751_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1751_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1751_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1751_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1763_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1763_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1763_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1763_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1763_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1775_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1775_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1775_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1775_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1775_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1801_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1801_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1801_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1801_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1801_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1957_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1957_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1957_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1957_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1957_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1986_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1986_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1986_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1986_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1986_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1986_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr57_1972 : std_logic_vector(31 downto 0);
    signal shr_1941 : std_logic_vector(31 downto 0);
    signal tmp10_1891 : std_logic_vector(15 downto 0);
    signal tmp113_1856 : std_logic_vector(15 downto 0);
    signal tmp114_1861 : std_logic_vector(15 downto 0);
    signal tmp115_1866 : std_logic_vector(15 downto 0);
    signal tmp11_1896 : std_logic_vector(15 downto 0);
    signal tmp12_1901 : std_logic_vector(15 downto 0);
    signal tmp14_1715 : std_logic_vector(15 downto 0);
    signal tmp17_1727 : std_logic_vector(15 downto 0);
    signal tmp1_1693 : std_logic_vector(15 downto 0);
    signal tmp20_1730 : std_logic_vector(15 downto 0);
    signal tmp26_1740 : std_logic_vector(15 downto 0);
    signal tmp29_1752 : std_logic_vector(15 downto 0);
    signal tmp2_1823 : std_logic_vector(15 downto 0);
    signal tmp39_1764 : std_logic_vector(15 downto 0);
    signal tmp3_1871 : std_logic_vector(15 downto 0);
    signal tmp43_1776 : std_logic_vector(15 downto 0);
    signal tmp4_1876 : std_logic_vector(15 downto 0);
    signal tmp54_1958 : std_logic_vector(63 downto 0);
    signal tmp5_1705 : std_logic_vector(15 downto 0);
    signal tmp6_1829 : std_logic_vector(15 downto 0);
    signal tmp7_1834 : std_logic_vector(15 downto 0);
    signal tmp83_1802 : std_logic_vector(15 downto 0);
    signal tmp8_1881 : std_logic_vector(15 downto 0);
    signal tmp9_1886 : std_logic_vector(15 downto 0);
    signal tmp_1818 : std_logic_vector(15 downto 0);
    signal type_cast_1788_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1810_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1816_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1827_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1841_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1843_wire : std_logic_vector(15 downto 0);
    signal type_cast_1848_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1850_wire : std_logic_vector(15 downto 0);
    signal type_cast_1907_wire : std_logic_vector(15 downto 0);
    signal type_cast_1910_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1915_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1930_wire : std_logic_vector(31 downto 0);
    signal type_cast_1935_wire : std_logic_vector(31 downto 0);
    signal type_cast_1938_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1945_wire : std_logic_vector(63 downto 0);
    signal type_cast_1961_wire : std_logic_vector(31 downto 0);
    signal type_cast_1966_wire : std_logic_vector(31 downto 0);
    signal type_cast_1969_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1975_wire : std_logic_vector(63 downto 0);
    signal type_cast_1991_wire : std_logic_vector(31 downto 0);
    signal type_cast_1997_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2002_wire : std_logic_vector(31 downto 0);
    signal type_cast_2004_wire : std_logic_vector(31 downto 0);
    signal type_cast_2017_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2025_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2030_wire : std_logic_vector(31 downto 0);
    signal type_cast_2050_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2056_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_1729_word_address_0 <= "0";
    array_obj_ref_1952_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1952_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1952_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1952_resized_base_address <= "00000000000000";
    array_obj_ref_1982_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1982_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1982_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1982_resized_base_address <= "00000000000000";
    iNsTr_10_1798 <= "00000000000000000000000000000100";
    iNsTr_2_1689 <= "00000000000000000000000000000110";
    iNsTr_3_1701 <= "00000000000000000000000000000101";
    iNsTr_4_1711 <= "00000000000000000000000000000000";
    iNsTr_5_1723 <= "00000000000000000000000000000101";
    iNsTr_6_1736 <= "00000000000000000000000000000001";
    iNsTr_7_1748 <= "00000000000000000000000000000110";
    iNsTr_8_1760 <= "00000000000000000000000000000110";
    iNsTr_9_1772 <= "00000000000000000000000000000101";
    ptr_deref_1692_word_offset_0 <= "0000000";
    ptr_deref_1704_word_offset_0 <= "0000000";
    ptr_deref_1714_word_offset_0 <= "0";
    ptr_deref_1726_word_offset_0 <= "0000000";
    ptr_deref_1739_word_offset_0 <= "0";
    ptr_deref_1751_word_offset_0 <= "0000000";
    ptr_deref_1763_word_offset_0 <= "0000000";
    ptr_deref_1775_word_offset_0 <= "0000000";
    ptr_deref_1801_word_offset_0 <= "0000000";
    ptr_deref_1957_word_offset_0 <= "00000000000000";
    ptr_deref_1986_word_offset_0 <= "00000000000000";
    type_cast_1788_wire_constant <= "00000000000000000000000000000001";
    type_cast_1810_wire_constant <= "00000000000000000000000000000001";
    type_cast_1816_wire_constant <= "1111111111111111";
    type_cast_1827_wire_constant <= "1111111111111111";
    type_cast_1841_wire_constant <= "0000000000000000";
    type_cast_1848_wire_constant <= "0000000000000000";
    type_cast_1910_wire_constant <= "0000000000000000";
    type_cast_1915_wire_constant <= "0000000000000100";
    type_cast_1938_wire_constant <= "00000000000000000000000000000010";
    type_cast_1969_wire_constant <= "00000000000000000000000000000010";
    type_cast_1997_wire_constant <= "00000000000000000000000000000100";
    type_cast_2017_wire_constant <= "0000000000000001";
    type_cast_2025_wire_constant <= "0000000000000001";
    type_cast_2050_wire_constant <= "0000000000000000";
    phi_stmt_1837: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1841_wire_constant & type_cast_1843_wire;
      req <= phi_stmt_1837_req_0 & phi_stmt_1837_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1837",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1837_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_1837,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1837
    phi_stmt_1844: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1848_wire_constant & type_cast_1850_wire;
      req <= phi_stmt_1844_req_0 & phi_stmt_1844_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1844",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1844_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_1844,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1844
    phi_stmt_1904: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1907_wire & type_cast_1910_wire_constant;
      req <= phi_stmt_1904_req_0 & phi_stmt_1904_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1904",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1904_ack_0,
          idata => idata,
          odata => indvar_1904,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1904
    -- flow-through select operator MUX_2052_inst
    input_dim1x_x2_2053 <= type_cast_2050_wire_constant when (cmp76_2037(0) /=  '0') else inc_2027;
    addr_of_1953_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1953_final_reg_req_0;
      addr_of_1953_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1953_final_reg_req_1;
      addr_of_1953_final_reg_ack_1<= rack(0);
      addr_of_1953_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1953_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1952_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1954,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1983_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1983_final_reg_req_0;
      addr_of_1983_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1983_final_reg_req_1;
      addr_of_1983_final_reg_ack_1<= rack(0);
      addr_of_1983_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1983_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1982_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx59_1984,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1779_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1779_inst_req_0;
      type_cast_1779_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1779_inst_req_1;
      type_cast_1779_inst_ack_1<= rack(0);
      type_cast_1779_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1779_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1_1693,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_1780,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1783_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1783_inst_req_0;
      type_cast_1783_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1783_inst_req_1;
      type_cast_1783_inst_ack_1<= rack(0);
      type_cast_1783_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1783_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp5_1705,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_1784,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1805_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1805_inst_req_0;
      type_cast_1805_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1805_inst_req_1;
      type_cast_1805_inst_ack_1<= rack(0);
      type_cast_1805_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1805_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp83_1802,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_1806,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1843_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1843_inst_req_0;
      type_cast_1843_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1843_inst_req_1;
      type_cast_1843_inst_ack_1<= rack(0);
      type_cast_1843_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1843_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2053,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1843_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1850_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1850_inst_req_0;
      type_cast_1850_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1850_inst_req_1;
      type_cast_1850_inst_ack_1<= rack(0);
      type_cast_1850_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1850_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc80x_xinput_dim0x_x2_2046,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1850_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1907_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1907_inst_req_0;
      type_cast_1907_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1907_inst_req_1;
      type_cast_1907_inst_ack_1<= rack(0);
      type_cast_1907_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1907_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2019,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1907_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1931_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1931_inst_req_0;
      type_cast_1931_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1931_inst_req_1;
      type_cast_1931_inst_ack_1<= rack(0);
      type_cast_1931_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1931_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1930_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_1932,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1935_inst
    process(conv53_1932) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv53_1932(31 downto 0);
      type_cast_1935_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1940_inst
    process(ASHR_i32_i32_1939_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1939_wire(31 downto 0);
      shr_1941 <= tmp_var; -- 
    end process;
    type_cast_1946_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1946_inst_req_0;
      type_cast_1946_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1946_inst_req_1;
      type_cast_1946_inst_ack_1<= rack(0);
      type_cast_1946_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1946_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1945_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1947,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1962_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1962_inst_req_0;
      type_cast_1962_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1962_inst_req_1;
      type_cast_1962_inst_ack_1<= rack(0);
      type_cast_1962_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1962_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1961_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_1963,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1966_inst
    process(conv56_1963) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv56_1963(31 downto 0);
      type_cast_1966_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1971_inst
    process(ASHR_i32_i32_1970_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1970_wire(31 downto 0);
      shr57_1972 <= tmp_var; -- 
    end process;
    type_cast_1976_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1976_inst_req_0;
      type_cast_1976_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1976_inst_req_1;
      type_cast_1976_inst_ack_1<= rack(0);
      type_cast_1976_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1976_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1975_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom58_1977,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1992_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1992_inst_req_0;
      type_cast_1992_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1992_inst_req_1;
      type_cast_1992_inst_ack_1<= rack(0);
      type_cast_1992_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1992_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1991_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_1993,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2002_inst
    process(add63_1999) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add63_1999(31 downto 0);
      type_cast_2002_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2004_inst
    process(conv65_1780) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv65_1780(31 downto 0);
      type_cast_2004_wire <= tmp_var; -- 
    end process;
    type_cast_2031_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2031_inst_req_0;
      type_cast_2031_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2031_inst_req_1;
      type_cast_2031_inst_ack_1<= rack(0);
      type_cast_2031_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2031_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2030_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2032,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2040_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2040_inst_req_0;
      type_cast_2040_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2040_inst_req_1;
      type_cast_2040_inst_ack_1<= rack(0);
      type_cast_2040_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2040_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp76_2037,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc80_2041,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2057_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2057_inst_req_0;
      type_cast_2057_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2057_inst_req_1;
      type_cast_2057_inst_ack_1<= rack(0);
      type_cast_2057_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2057_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2056_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_2058,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_1729_gather_scatter
    process(LOAD_padding_1729_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_1729_data_0;
      ov(15 downto 0) := iv;
      tmp20_1730 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1952_index_1_rename
    process(R_idxprom_1951_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1951_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1951_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1952_index_1_resize
    process(idxprom_1947) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1947;
      ov := iv(13 downto 0);
      R_idxprom_1951_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1952_root_address_inst
    process(array_obj_ref_1952_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1952_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1952_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1982_index_1_rename
    process(R_idxprom58_1981_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom58_1981_resized;
      ov(13 downto 0) := iv;
      R_idxprom58_1981_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1982_index_1_resize
    process(idxprom58_1977) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom58_1977;
      ov := iv(13 downto 0);
      R_idxprom58_1981_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1982_root_address_inst
    process(array_obj_ref_1982_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1982_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1982_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1692_addr_0
    process(ptr_deref_1692_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1692_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1692_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1692_base_resize
    process(iNsTr_2_1689) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1689;
      ov := iv(6 downto 0);
      ptr_deref_1692_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1692_gather_scatter
    process(ptr_deref_1692_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1692_data_0;
      ov(15 downto 0) := iv;
      tmp1_1693 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1692_root_address_inst
    process(ptr_deref_1692_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1692_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1692_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1704_addr_0
    process(ptr_deref_1704_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1704_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1704_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1704_base_resize
    process(iNsTr_3_1701) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_1701;
      ov := iv(6 downto 0);
      ptr_deref_1704_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1704_gather_scatter
    process(ptr_deref_1704_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1704_data_0;
      ov(15 downto 0) := iv;
      tmp5_1705 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1704_root_address_inst
    process(ptr_deref_1704_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1704_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1704_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1714_addr_0
    process(ptr_deref_1714_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1714_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1714_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1714_base_resize
    process(iNsTr_4_1711) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_1711;
      ov := iv(0 downto 0);
      ptr_deref_1714_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1714_gather_scatter
    process(ptr_deref_1714_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1714_data_0;
      ov(15 downto 0) := iv;
      tmp14_1715 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1714_root_address_inst
    process(ptr_deref_1714_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1714_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1714_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1726_addr_0
    process(ptr_deref_1726_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1726_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1726_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1726_base_resize
    process(iNsTr_5_1723) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_1723;
      ov := iv(6 downto 0);
      ptr_deref_1726_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1726_gather_scatter
    process(ptr_deref_1726_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1726_data_0;
      ov(15 downto 0) := iv;
      tmp17_1727 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1726_root_address_inst
    process(ptr_deref_1726_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1726_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1726_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1739_addr_0
    process(ptr_deref_1739_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1739_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1739_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1739_base_resize
    process(iNsTr_6_1736) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_1736;
      ov := iv(0 downto 0);
      ptr_deref_1739_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1739_gather_scatter
    process(ptr_deref_1739_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1739_data_0;
      ov(15 downto 0) := iv;
      tmp26_1740 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1739_root_address_inst
    process(ptr_deref_1739_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1739_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1739_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1751_addr_0
    process(ptr_deref_1751_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1751_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1751_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1751_base_resize
    process(iNsTr_7_1748) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_1748;
      ov := iv(6 downto 0);
      ptr_deref_1751_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1751_gather_scatter
    process(ptr_deref_1751_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1751_data_0;
      ov(15 downto 0) := iv;
      tmp29_1752 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1751_root_address_inst
    process(ptr_deref_1751_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1751_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1751_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1763_addr_0
    process(ptr_deref_1763_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1763_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1763_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1763_base_resize
    process(iNsTr_8_1760) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_1760;
      ov := iv(6 downto 0);
      ptr_deref_1763_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1763_gather_scatter
    process(ptr_deref_1763_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1763_data_0;
      ov(15 downto 0) := iv;
      tmp39_1764 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1763_root_address_inst
    process(ptr_deref_1763_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1763_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1763_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1775_addr_0
    process(ptr_deref_1775_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1775_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1775_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1775_base_resize
    process(iNsTr_9_1772) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_1772;
      ov := iv(6 downto 0);
      ptr_deref_1775_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1775_gather_scatter
    process(ptr_deref_1775_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1775_data_0;
      ov(15 downto 0) := iv;
      tmp43_1776 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1775_root_address_inst
    process(ptr_deref_1775_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1775_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1775_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1801_addr_0
    process(ptr_deref_1801_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1801_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1801_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1801_base_resize
    process(iNsTr_10_1798) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_1798;
      ov := iv(6 downto 0);
      ptr_deref_1801_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1801_gather_scatter
    process(ptr_deref_1801_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1801_data_0;
      ov(15 downto 0) := iv;
      tmp83_1802 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1801_root_address_inst
    process(ptr_deref_1801_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1801_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1801_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1957_addr_0
    process(ptr_deref_1957_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1957_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1957_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1957_base_resize
    process(arrayidx_1954) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1954;
      ov := iv(13 downto 0);
      ptr_deref_1957_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1957_gather_scatter
    process(ptr_deref_1957_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1957_data_0;
      ov(63 downto 0) := iv;
      tmp54_1958 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1957_root_address_inst
    process(ptr_deref_1957_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1957_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1957_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1986_addr_0
    process(ptr_deref_1986_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1986_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1986_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1986_base_resize
    process(arrayidx59_1984) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx59_1984;
      ov := iv(13 downto 0);
      ptr_deref_1986_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1986_gather_scatter
    process(tmp54_1958) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp54_1958;
      ov(63 downto 0) := iv;
      ptr_deref_1986_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1986_root_address_inst
    process(ptr_deref_1986_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1986_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1986_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2007_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2006;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2007_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2007_branch_req_0,
          ack0 => if_stmt_2007_branch_ack_0,
          ack1 => if_stmt_2007_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2064_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp86_2063;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2064_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2064_branch_req_0,
          ack0 => if_stmt_2064_branch_ack_0,
          ack1 => if_stmt_2064_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1817_inst
    process(tmp29_1752) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp29_1752, type_cast_1816_wire_constant, tmp_var);
      tmp_1818 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1828_inst
    process(tmp17_1727) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp17_1727, type_cast_1827_wire_constant, tmp_var);
      tmp6_1829 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1860_inst
    process(input_dim1x_x1x_xph_1837, tmp113_1856) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1837, tmp113_1856, tmp_var);
      tmp114_1861 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1875_inst
    process(tmp2_1823, tmp3_1871) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp2_1823, tmp3_1871, tmp_var);
      tmp4_1876 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1885_inst
    process(tmp7_1834, tmp8_1881) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp7_1834, tmp8_1881, tmp_var);
      tmp9_1886 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1895_inst
    process(tmp4_1876, tmp10_1891) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp4_1876, tmp10_1891, tmp_var);
      tmp11_1896 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1921_inst
    process(tmp115_1866, input_dim2x_x1_1917) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp115_1866, input_dim2x_x1_1917, tmp_var);
      add10_1922 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1926_inst
    process(tmp12_1901, input_dim2x_x1_1917) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp12_1901, input_dim2x_x1_1917, tmp_var);
      add50_1927 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2018_inst
    process(indvar_1904) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1904, type_cast_2017_wire_constant, tmp_var);
      indvarx_xnext_2019 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2026_inst
    process(input_dim1x_x1x_xph_1837) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1837, type_cast_2025_wire_constant, tmp_var);
      inc_2027 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2045_inst
    process(inc80_2041, input_dim0x_x2x_xph_1844) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc80_2041, input_dim0x_x2x_xph_1844, tmp_var);
      inc80x_xinput_dim0x_x2_2046 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1998_inst
    process(conv62_1993) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv62_1993, type_cast_1997_wire_constant, tmp_var);
      add63_1999 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1939_inst
    process(type_cast_1935_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1935_wire, type_cast_1938_wire_constant, tmp_var);
      ASHR_i32_i32_1939_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1970_inst
    process(type_cast_1966_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1966_wire, type_cast_1969_wire_constant, tmp_var);
      ASHR_i32_i32_1970_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2036_inst
    process(conv73_2032, div_1790) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv73_2032, div_1790, tmp_var);
      cmp76_2037 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2062_inst
    process(conv82_2058, div85_1812) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv82_2058, div85_1812, tmp_var);
      cmp86_2063 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1789_inst
    process(conv75_1784) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv75_1784, type_cast_1788_wire_constant, tmp_var);
      div_1790 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1811_inst
    process(conv84_1806) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv84_1806, type_cast_1810_wire_constant, tmp_var);
      div85_1812 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1855_inst
    process(tmp5_1705, input_dim0x_x2x_xph_1844) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp5_1705, input_dim0x_x2x_xph_1844, tmp_var);
      tmp113_1856 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1865_inst
    process(tmp1_1693, tmp114_1861) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_1693, tmp114_1861, tmp_var);
      tmp115_1866 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1870_inst
    process(tmp26_1740, input_dim1x_x1x_xph_1837) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp26_1740, input_dim1x_x1x_xph_1837, tmp_var);
      tmp3_1871 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1880_inst
    process(tmp14_1715, input_dim0x_x2x_xph_1844) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp14_1715, input_dim0x_x2x_xph_1844, tmp_var);
      tmp8_1881 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1890_inst
    process(tmp43_1776, tmp9_1886) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp43_1776, tmp9_1886, tmp_var);
      tmp10_1891 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1900_inst
    process(tmp39_1764, tmp11_1896) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp39_1764, tmp11_1896, tmp_var);
      tmp12_1901 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1916_inst
    process(indvar_1904) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1904, type_cast_1915_wire_constant, tmp_var);
      input_dim2x_x1_1917 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2005_inst
    process(type_cast_2002_wire, type_cast_2004_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2002_wire, type_cast_2004_wire, tmp_var);
      cmp_2006 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1822_inst
    process(tmp_1818, tmp20_1730) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp_1818, tmp20_1730, tmp_var);
      tmp2_1823 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1833_inst
    process(tmp6_1829, tmp20_1730) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp6_1829, tmp20_1730, tmp_var);
      tmp7_1834 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_1952_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1951_scaled;
      array_obj_ref_1952_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1952_index_offset_req_0;
      array_obj_ref_1952_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1952_index_offset_req_1;
      array_obj_ref_1952_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_1982_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom58_1981_scaled;
      array_obj_ref_1982_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1982_index_offset_req_0;
      array_obj_ref_1982_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1982_index_offset_req_1;
      array_obj_ref_1982_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- unary operator type_cast_1930_inst
    process(add10_1922) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add10_1922, tmp_var);
      type_cast_1930_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1945_inst
    process(shr_1941) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1941, tmp_var);
      type_cast_1945_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1961_inst
    process(add50_1927) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add50_1927, tmp_var);
      type_cast_1961_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1975_inst
    process(shr57_1972) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr57_1972, tmp_var);
      type_cast_1975_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1991_inst
    process(input_dim2x_x1_1917) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_1917, tmp_var);
      type_cast_1991_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2030_inst
    process(inc_2027) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2027, tmp_var);
      type_cast_2030_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2056_inst
    process(inc80x_xinput_dim0x_x2_2046) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc80x_xinput_dim0x_x2_2046, tmp_var);
      type_cast_2056_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_1729_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_1729_load_0_req_0;
      LOAD_padding_1729_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_1729_load_0_req_1;
      LOAD_padding_1729_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_1729_word_address_0;
      LOAD_padding_1729_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1692_load_0 ptr_deref_1704_load_0 ptr_deref_1801_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1692_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1704_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1801_load_0_req_0;
      ptr_deref_1692_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1704_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1801_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1692_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1704_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1801_load_0_req_1;
      ptr_deref_1692_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1704_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1801_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1692_word_address_0 & ptr_deref_1704_word_address_0 & ptr_deref_1801_word_address_0;
      ptr_deref_1692_data_0 <= data_out(47 downto 32);
      ptr_deref_1704_data_0 <= data_out(31 downto 16);
      ptr_deref_1801_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 16,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(15 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_1714_load_0 ptr_deref_1739_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1714_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1739_load_0_req_0;
      ptr_deref_1714_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1739_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1714_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1739_load_0_req_1;
      ptr_deref_1714_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1739_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1714_word_address_0 & ptr_deref_1739_word_address_0;
      ptr_deref_1714_data_0 <= data_out(31 downto 16);
      ptr_deref_1739_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(15 downto 0),
          mtag => memory_space_8_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_1726_load_0 ptr_deref_1751_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1726_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1751_load_0_req_0;
      ptr_deref_1726_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1751_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1726_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1751_load_0_req_1;
      ptr_deref_1726_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1751_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1726_word_address_0 & ptr_deref_1751_word_address_0;
      ptr_deref_1726_data_0 <= data_out(31 downto 16);
      ptr_deref_1751_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(15 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_1763_load_0 ptr_deref_1775_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1763_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1775_load_0_req_0;
      ptr_deref_1763_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1775_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1763_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1775_load_0_req_1;
      ptr_deref_1763_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1775_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1763_word_address_0 & ptr_deref_1775_word_address_0;
      ptr_deref_1763_data_0 <= data_out(31 downto 16);
      ptr_deref_1775_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(15 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_1957_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1957_load_0_req_0;
      ptr_deref_1957_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1957_load_0_req_1;
      ptr_deref_1957_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1957_word_address_0;
      ptr_deref_1957_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(13 downto 0),
          mtag => memory_space_4_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(63 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_1986_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1986_store_0_req_0;
      ptr_deref_1986_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1986_store_0_req_1;
      ptr_deref_1986_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1986_word_address_0;
      data_in <= ptr_deref_1986_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(13 downto 0),
          mdata => memory_space_6_sr_data(63 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1679_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_start_1679_inst_req_0;
      RPIPE_Block0_start_1679_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_start_1679_inst_req_1;
      RPIPE_Block0_start_1679_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_1680 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_2072_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_2072_inst_req_0;
      WPIPE_Block0_done_2072_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_2072_inst_req_1;
      WPIPE_Block0_done_2072_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1680;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_6188_start: Boolean;
  signal convTransposeB_CP_6188_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_2148_load_0_ack_0 : boolean;
  signal ptr_deref_2148_load_0_req_1 : boolean;
  signal ptr_deref_2148_load_0_ack_1 : boolean;
  signal ptr_deref_2160_load_0_req_0 : boolean;
  signal ptr_deref_2160_load_0_ack_0 : boolean;
  signal type_cast_2192_inst_ack_1 : boolean;
  signal type_cast_2188_inst_req_0 : boolean;
  signal type_cast_2188_inst_ack_0 : boolean;
  signal ptr_deref_2184_load_0_req_0 : boolean;
  signal ptr_deref_2184_load_0_ack_0 : boolean;
  signal type_cast_2188_inst_req_1 : boolean;
  signal type_cast_2188_inst_ack_1 : boolean;
  signal ptr_deref_2172_load_0_req_1 : boolean;
  signal type_cast_2192_inst_req_0 : boolean;
  signal type_cast_2192_inst_ack_0 : boolean;
  signal type_cast_2192_inst_req_1 : boolean;
  signal ptr_deref_2172_load_0_ack_1 : boolean;
  signal ptr_deref_2160_load_0_req_1 : boolean;
  signal ptr_deref_2160_load_0_ack_1 : boolean;
  signal ptr_deref_2148_load_0_req_0 : boolean;
  signal ptr_deref_2184_load_0_req_1 : boolean;
  signal ptr_deref_2184_load_0_ack_1 : boolean;
  signal ptr_deref_2204_load_0_req_1 : boolean;
  signal ptr_deref_2204_load_0_ack_1 : boolean;
  signal ptr_deref_2204_load_0_req_0 : boolean;
  signal ptr_deref_2204_load_0_ack_0 : boolean;
  signal ptr_deref_2172_load_0_ack_0 : boolean;
  signal ptr_deref_2172_load_0_req_0 : boolean;
  signal RPIPE_Block1_start_2082_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2082_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2082_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2082_inst_ack_1 : boolean;
  signal ptr_deref_2095_load_0_req_0 : boolean;
  signal ptr_deref_2095_load_0_ack_0 : boolean;
  signal ptr_deref_2095_load_0_req_1 : boolean;
  signal ptr_deref_2095_load_0_ack_1 : boolean;
  signal ptr_deref_2113_load_0_req_0 : boolean;
  signal ptr_deref_2113_load_0_ack_0 : boolean;
  signal ptr_deref_2113_load_0_req_1 : boolean;
  signal ptr_deref_2113_load_0_ack_1 : boolean;
  signal ptr_deref_2123_load_0_req_0 : boolean;
  signal ptr_deref_2123_load_0_ack_0 : boolean;
  signal ptr_deref_2123_load_0_req_1 : boolean;
  signal ptr_deref_2123_load_0_ack_1 : boolean;
  signal ptr_deref_2135_load_0_req_0 : boolean;
  signal ptr_deref_2135_load_0_ack_0 : boolean;
  signal ptr_deref_2135_load_0_req_1 : boolean;
  signal ptr_deref_2135_load_0_ack_1 : boolean;
  signal LOAD_padding_2138_load_0_req_0 : boolean;
  signal LOAD_padding_2138_load_0_ack_0 : boolean;
  signal LOAD_padding_2138_load_0_req_1 : boolean;
  signal LOAD_padding_2138_load_0_ack_1 : boolean;
  signal type_cast_2208_inst_req_0 : boolean;
  signal type_cast_2208_inst_ack_0 : boolean;
  signal type_cast_2208_inst_req_1 : boolean;
  signal type_cast_2208_inst_ack_1 : boolean;
  signal type_cast_2333_inst_req_0 : boolean;
  signal type_cast_2333_inst_ack_0 : boolean;
  signal type_cast_2333_inst_req_1 : boolean;
  signal type_cast_2333_inst_ack_1 : boolean;
  signal type_cast_2347_inst_req_0 : boolean;
  signal type_cast_2347_inst_ack_0 : boolean;
  signal type_cast_2347_inst_req_1 : boolean;
  signal type_cast_2347_inst_ack_1 : boolean;
  signal array_obj_ref_2353_index_offset_req_0 : boolean;
  signal array_obj_ref_2353_index_offset_ack_0 : boolean;
  signal array_obj_ref_2353_index_offset_req_1 : boolean;
  signal array_obj_ref_2353_index_offset_ack_1 : boolean;
  signal addr_of_2354_final_reg_req_0 : boolean;
  signal addr_of_2354_final_reg_ack_0 : boolean;
  signal addr_of_2354_final_reg_req_1 : boolean;
  signal addr_of_2354_final_reg_ack_1 : boolean;
  signal ptr_deref_2358_load_0_req_0 : boolean;
  signal ptr_deref_2358_load_0_ack_0 : boolean;
  signal ptr_deref_2358_load_0_req_1 : boolean;
  signal ptr_deref_2358_load_0_ack_1 : boolean;
  signal type_cast_2363_inst_req_0 : boolean;
  signal type_cast_2363_inst_ack_0 : boolean;
  signal type_cast_2363_inst_req_1 : boolean;
  signal type_cast_2363_inst_ack_1 : boolean;
  signal type_cast_2377_inst_req_0 : boolean;
  signal type_cast_2377_inst_ack_0 : boolean;
  signal type_cast_2377_inst_req_1 : boolean;
  signal type_cast_2377_inst_ack_1 : boolean;
  signal array_obj_ref_2383_index_offset_req_0 : boolean;
  signal array_obj_ref_2383_index_offset_ack_0 : boolean;
  signal array_obj_ref_2383_index_offset_req_1 : boolean;
  signal array_obj_ref_2383_index_offset_ack_1 : boolean;
  signal addr_of_2384_final_reg_req_0 : boolean;
  signal addr_of_2384_final_reg_ack_0 : boolean;
  signal addr_of_2384_final_reg_req_1 : boolean;
  signal addr_of_2384_final_reg_ack_1 : boolean;
  signal ptr_deref_2387_store_0_req_0 : boolean;
  signal ptr_deref_2387_store_0_ack_0 : boolean;
  signal ptr_deref_2387_store_0_req_1 : boolean;
  signal ptr_deref_2387_store_0_ack_1 : boolean;
  signal type_cast_2393_inst_req_0 : boolean;
  signal type_cast_2393_inst_ack_0 : boolean;
  signal type_cast_2393_inst_req_1 : boolean;
  signal type_cast_2393_inst_ack_1 : boolean;
  signal if_stmt_2408_branch_req_0 : boolean;
  signal if_stmt_2408_branch_ack_1 : boolean;
  signal if_stmt_2408_branch_ack_0 : boolean;
  signal type_cast_2432_inst_req_0 : boolean;
  signal type_cast_2432_inst_ack_0 : boolean;
  signal type_cast_2432_inst_req_1 : boolean;
  signal type_cast_2432_inst_ack_1 : boolean;
  signal type_cast_2466_inst_req_0 : boolean;
  signal type_cast_2466_inst_ack_0 : boolean;
  signal type_cast_2466_inst_req_1 : boolean;
  signal type_cast_2466_inst_ack_1 : boolean;
  signal if_stmt_2473_branch_req_0 : boolean;
  signal if_stmt_2473_branch_ack_1 : boolean;
  signal if_stmt_2473_branch_ack_0 : boolean;
  signal WPIPE_Block1_done_2481_inst_req_0 : boolean;
  signal WPIPE_Block1_done_2481_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_2481_inst_req_1 : boolean;
  signal WPIPE_Block1_done_2481_inst_ack_1 : boolean;
  signal type_cast_2243_inst_req_0 : boolean;
  signal type_cast_2243_inst_ack_0 : boolean;
  signal type_cast_2243_inst_req_1 : boolean;
  signal type_cast_2243_inst_ack_1 : boolean;
  signal phi_stmt_2240_req_0 : boolean;
  signal phi_stmt_2246_req_0 : boolean;
  signal type_cast_2245_inst_req_0 : boolean;
  signal type_cast_2245_inst_ack_0 : boolean;
  signal type_cast_2245_inst_req_1 : boolean;
  signal type_cast_2245_inst_ack_1 : boolean;
  signal phi_stmt_2240_req_1 : boolean;
  signal type_cast_2252_inst_req_0 : boolean;
  signal type_cast_2252_inst_ack_0 : boolean;
  signal type_cast_2252_inst_req_1 : boolean;
  signal type_cast_2252_inst_ack_1 : boolean;
  signal phi_stmt_2246_req_1 : boolean;
  signal phi_stmt_2240_ack_0 : boolean;
  signal phi_stmt_2246_ack_0 : boolean;
  signal type_cast_2309_inst_req_0 : boolean;
  signal type_cast_2309_inst_ack_0 : boolean;
  signal type_cast_2309_inst_req_1 : boolean;
  signal type_cast_2309_inst_ack_1 : boolean;
  signal phi_stmt_2306_req_0 : boolean;
  signal phi_stmt_2306_req_1 : boolean;
  signal phi_stmt_2306_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_6188_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_6188_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_6188_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_6188_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_6188: Block -- control-path 
    signal convTransposeB_CP_6188_elements: BooleanArray(85 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_6188_elements(0) <= convTransposeB_CP_6188_start;
    convTransposeB_CP_6188_symbol <= convTransposeB_CP_6188_elements(63);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2080/$entry
      -- CP-element group 0: 	 branch_block_stmt_2080/branch_block_stmt_2080__entry__
      -- CP-element group 0: 	 branch_block_stmt_2080/assign_stmt_2083__entry__
      -- CP-element group 0: 	 branch_block_stmt_2080/assign_stmt_2083/$entry
      -- CP-element group 0: 	 branch_block_stmt_2080/assign_stmt_2083/RPIPE_Block1_start_2082_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2080/assign_stmt_2083/RPIPE_Block1_start_2082_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2080/assign_stmt_2083/RPIPE_Block1_start_2082_Sample/rr
      -- 
    rr_6236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(0), ack => RPIPE_Block1_start_2082_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2080/assign_stmt_2083/RPIPE_Block1_start_2082_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_2080/assign_stmt_2083/RPIPE_Block1_start_2082_update_start_
      -- CP-element group 1: 	 branch_block_stmt_2080/assign_stmt_2083/RPIPE_Block1_start_2082_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_2080/assign_stmt_2083/RPIPE_Block1_start_2082_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_2080/assign_stmt_2083/RPIPE_Block1_start_2082_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2080/assign_stmt_2083/RPIPE_Block1_start_2082_Update/cr
      -- 
    ra_6237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2082_inst_ack_0, ack => convTransposeB_CP_6188_elements(1)); -- 
    cr_6241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(1), ack => RPIPE_Block1_start_2082_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	25 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2:  members (262) 
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2188_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2188_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2192_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2192_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2188_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2192_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2083__exit__
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237__entry__
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2083/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2083/RPIPE_Block1_start_2082_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2083/RPIPE_Block1_start_2082_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2083/RPIPE_Block1_start_2082_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2208_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2208_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2208_Update/cr
      -- 
    ca_6242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2082_inst_ack_1, ack => convTransposeB_CP_6188_elements(2)); -- 
    cr_6522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => ptr_deref_2148_load_0_req_1); -- 
    rr_6561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => ptr_deref_2160_load_0_req_0); -- 
    rr_6661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => ptr_deref_2184_load_0_req_0); -- 
    cr_6691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => type_cast_2188_inst_req_1); -- 
    cr_6622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => ptr_deref_2172_load_0_req_1); -- 
    cr_6705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => type_cast_2192_inst_req_1); -- 
    cr_6572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => ptr_deref_2160_load_0_req_1); -- 
    rr_6511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => ptr_deref_2148_load_0_req_0); -- 
    cr_6672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => ptr_deref_2184_load_0_req_1); -- 
    cr_6750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => ptr_deref_2204_load_0_req_1); -- 
    rr_6739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => ptr_deref_2204_load_0_req_0); -- 
    rr_6611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => ptr_deref_2172_load_0_req_0); -- 
    rr_6278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => ptr_deref_2095_load_0_req_0); -- 
    cr_6289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => ptr_deref_2095_load_0_req_1); -- 
    rr_6328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => ptr_deref_2113_load_0_req_0); -- 
    cr_6339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => ptr_deref_2113_load_0_req_1); -- 
    rr_6378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => ptr_deref_2123_load_0_req_0); -- 
    cr_6389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => ptr_deref_2123_load_0_req_1); -- 
    rr_6428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => ptr_deref_2135_load_0_req_0); -- 
    cr_6439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => ptr_deref_2135_load_0_req_1); -- 
    rr_6461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => LOAD_padding_2138_load_0_req_0); -- 
    cr_6472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => LOAD_padding_2138_load_0_req_1); -- 
    cr_6769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(2), ack => type_cast_2208_inst_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_Sample/word_access_start/word_0/ra
      -- 
    ra_6279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2095_load_0_ack_0, ack => convTransposeB_CP_6188_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	23 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2192_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2192_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2192_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_Update/ptr_deref_2095_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_Update/ptr_deref_2095_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_Update/ptr_deref_2095_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2095_Update/ptr_deref_2095_Merge/merge_ack
      -- 
    ca_6290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2095_load_0_ack_1, ack => convTransposeB_CP_6188_elements(4)); -- 
    rr_6700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(4), ack => type_cast_2192_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_Sample/word_access_start/word_0/ra
      -- 
    ra_6329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2113_load_0_ack_0, ack => convTransposeB_CP_6188_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	21 
    -- CP-element group 6:  members (12) 
      -- CP-element group 6: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2188_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2188_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2188_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_Update/ptr_deref_2113_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_Update/ptr_deref_2113_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_Update/ptr_deref_2113_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2113_Update/ptr_deref_2113_Merge/merge_ack
      -- 
    ca_6340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2113_load_0_ack_1, ack => convTransposeB_CP_6188_elements(6)); -- 
    rr_6686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(6), ack => type_cast_2188_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_Sample/word_access_start/word_0/ra
      -- 
    ra_6379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2123_load_0_ack_0, ack => convTransposeB_CP_6188_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	29 
    -- CP-element group 8:  members (9) 
      -- CP-element group 8: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_Update/ptr_deref_2123_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_Update/ptr_deref_2123_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_Update/ptr_deref_2123_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2123_Update/ptr_deref_2123_Merge/merge_ack
      -- 
    ca_6390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2123_load_0_ack_1, ack => convTransposeB_CP_6188_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_Sample/word_access_start/word_0/ra
      -- 
    ra_6429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2135_load_0_ack_0, ack => convTransposeB_CP_6188_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	29 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_Update/ptr_deref_2135_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_Update/ptr_deref_2135_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_Update/ptr_deref_2135_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2135_Update/ptr_deref_2135_Merge/merge_ack
      -- 
    ca_6440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2135_load_0_ack_1, ack => convTransposeB_CP_6188_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_Sample/word_access_start/word_0/ra
      -- 
    ra_6462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2138_load_0_ack_0, ack => convTransposeB_CP_6188_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	29 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_Update/LOAD_padding_2138_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_Update/LOAD_padding_2138_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_Update/LOAD_padding_2138_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/LOAD_padding_2138_Update/LOAD_padding_2138_Merge/merge_ack
      -- 
    ca_6473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2138_load_0_ack_1, ack => convTransposeB_CP_6188_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_Sample/word_access_start/word_0/ra
      -- CP-element group 13: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_sample_completed_
      -- 
    ra_6512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2148_load_0_ack_0, ack => convTransposeB_CP_6188_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	29 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_Update/ptr_deref_2148_Merge/merge_ack
      -- CP-element group 14: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_Update/ptr_deref_2148_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_Update/ptr_deref_2148_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_Update/ptr_deref_2148_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2148_update_completed_
      -- 
    ca_6523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2148_load_0_ack_1, ack => convTransposeB_CP_6188_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_Sample/word_access_start/word_0/ra
      -- 
    ra_6562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2160_load_0_ack_0, ack => convTransposeB_CP_6188_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	29 
    -- CP-element group 16:  members (9) 
      -- CP-element group 16: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_Update/ptr_deref_2160_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_Update/ptr_deref_2160_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_Update/ptr_deref_2160_Merge/merge_ack
      -- CP-element group 16: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2160_Update/ptr_deref_2160_Merge/merge_req
      -- 
    ca_6573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2160_load_0_ack_1, ack => convTransposeB_CP_6188_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_Sample/word_access_start/word_0/ra
      -- 
    ra_6612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2172_load_0_ack_0, ack => convTransposeB_CP_6188_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	29 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_Update/ptr_deref_2172_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_Update/ptr_deref_2172_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_Update/ptr_deref_2172_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2172_Update/ptr_deref_2172_Merge/merge_ack
      -- 
    ca_6623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2172_load_0_ack_1, ack => convTransposeB_CP_6188_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_Sample/word_access_start/word_0/ra
      -- CP-element group 19: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_sample_completed_
      -- 
    ra_6662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2184_load_0_ack_0, ack => convTransposeB_CP_6188_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	29 
    -- CP-element group 20:  members (9) 
      -- CP-element group 20: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_Update/ptr_deref_2184_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_Update/ptr_deref_2184_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_Update/ptr_deref_2184_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_Update/ptr_deref_2184_Merge/merge_ack
      -- CP-element group 20: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2184_Update/word_access_complete/word_0/ca
      -- 
    ca_6673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2184_load_0_ack_1, ack => convTransposeB_CP_6188_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	6 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2188_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2188_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2188_sample_completed_
      -- 
    ra_6687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2188_inst_ack_0, ack => convTransposeB_CP_6188_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	29 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2188_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2188_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2188_Update/$exit
      -- 
    ca_6692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2188_inst_ack_1, ack => convTransposeB_CP_6188_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	4 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2192_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2192_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2192_sample_completed_
      -- 
    ra_6701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2192_inst_ack_0, ack => convTransposeB_CP_6188_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	29 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2192_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2192_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2192_Update/$exit
      -- 
    ca_6706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2192_inst_ack_1, ack => convTransposeB_CP_6188_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_Sample/word_access_start/word_0/ra
      -- 
    ra_6740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2204_load_0_ack_0, ack => convTransposeB_CP_6188_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (12) 
      -- CP-element group 26: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_Update/word_access_complete/word_0/ca
      -- CP-element group 26: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_Update/ptr_deref_2204_Merge/$entry
      -- CP-element group 26: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_Update/ptr_deref_2204_Merge/$exit
      -- CP-element group 26: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_Update/ptr_deref_2204_Merge/merge_req
      -- CP-element group 26: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_Update/ptr_deref_2204_Merge/merge_ack
      -- CP-element group 26: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/ptr_deref_2204_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2208_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2208_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2208_Sample/rr
      -- 
    ca_6751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2204_load_0_ack_1, ack => convTransposeB_CP_6188_elements(26)); -- 
    rr_6764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(26), ack => type_cast_2208_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2208_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2208_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2208_Sample/ra
      -- 
    ra_6765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2208_inst_ack_0, ack => convTransposeB_CP_6188_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2208_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2208_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/type_cast_2208_Update/ca
      -- 
    ca_6770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2208_inst_ack_1, ack => convTransposeB_CP_6188_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  place  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	18 
    -- CP-element group 29: 	22 
    -- CP-element group 29: 	16 
    -- CP-element group 29: 	8 
    -- CP-element group 29: 	28 
    -- CP-element group 29: 	20 
    -- CP-element group 29: 	24 
    -- CP-element group 29: 	10 
    -- CP-element group 29: 	12 
    -- CP-element group 29: 	14 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	65 
    -- CP-element group 29: 	67 
    -- CP-element group 29: 	64 
    -- CP-element group 29:  members (14) 
      -- CP-element group 29: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237__exit__
      -- CP-element group 29: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter
      -- CP-element group 29: 	 branch_block_stmt_2080/assign_stmt_2092_to_assign_stmt_2237/$exit
      -- CP-element group 29: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 29: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/$entry
      -- CP-element group 29: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/$entry
      -- CP-element group 29: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/SplitProtocol/$entry
      -- CP-element group 29: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/SplitProtocol/Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/SplitProtocol/Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/SplitProtocol/Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/SplitProtocol/Update/cr
      -- CP-element group 29: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/$entry
      -- CP-element group 29: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/phi_stmt_2246_sources/$entry
      -- 
    rr_7146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(29), ack => type_cast_2243_inst_req_0); -- 
    cr_7151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(29), ack => type_cast_2243_inst_req_1); -- 
    convTransposeB_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeB_CP_6188_elements(18) & convTransposeB_CP_6188_elements(22) & convTransposeB_CP_6188_elements(16) & convTransposeB_CP_6188_elements(8) & convTransposeB_CP_6188_elements(28) & convTransposeB_CP_6188_elements(20) & convTransposeB_CP_6188_elements(24) & convTransposeB_CP_6188_elements(10) & convTransposeB_CP_6188_elements(12) & convTransposeB_CP_6188_elements(14);
      gj_convTransposeB_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_6188_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	85 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2333_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2333_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2333_Sample/ra
      -- 
    ra_6785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2333_inst_ack_0, ack => convTransposeB_CP_6188_elements(30)); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	85 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2333_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2333_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2333_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2347_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2347_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2347_Sample/rr
      -- 
    ca_6790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2333_inst_ack_1, ack => convTransposeB_CP_6188_elements(31)); -- 
    rr_6798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(31), ack => type_cast_2347_inst_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2347_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2347_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2347_Sample/ra
      -- 
    ra_6799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2347_inst_ack_0, ack => convTransposeB_CP_6188_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	85 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (16) 
      -- CP-element group 33: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2347_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2347_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2347_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_index_resized_1
      -- CP-element group 33: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_index_scaled_1
      -- CP-element group 33: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_index_computed_1
      -- CP-element group 33: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_index_resize_1/$entry
      -- CP-element group 33: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_index_resize_1/$exit
      -- CP-element group 33: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_index_resize_1/index_resize_req
      -- CP-element group 33: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_index_resize_1/index_resize_ack
      -- CP-element group 33: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_index_scale_1/$entry
      -- CP-element group 33: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_index_scale_1/$exit
      -- CP-element group 33: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_index_scale_1/scale_rename_req
      -- CP-element group 33: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_index_scale_1/scale_rename_ack
      -- CP-element group 33: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_final_index_sum_regn_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_final_index_sum_regn_Sample/req
      -- 
    ca_6804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2347_inst_ack_1, ack => convTransposeB_CP_6188_elements(33)); -- 
    req_6829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(33), ack => array_obj_ref_2353_index_offset_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	53 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_final_index_sum_regn_sample_complete
      -- CP-element group 34: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_final_index_sum_regn_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_final_index_sum_regn_Sample/ack
      -- 
    ack_6830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2353_index_offset_ack_0, ack => convTransposeB_CP_6188_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	85 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (11) 
      -- CP-element group 35: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2354_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_root_address_calculated
      -- CP-element group 35: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_offset_calculated
      -- CP-element group 35: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_final_index_sum_regn_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_final_index_sum_regn_Update/ack
      -- CP-element group 35: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_base_plus_offset/$entry
      -- CP-element group 35: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_base_plus_offset/$exit
      -- CP-element group 35: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_base_plus_offset/sum_rename_req
      -- CP-element group 35: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_base_plus_offset/sum_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2354_request/$entry
      -- CP-element group 35: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2354_request/req
      -- 
    ack_6835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2353_index_offset_ack_1, ack => convTransposeB_CP_6188_elements(35)); -- 
    req_6844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(35), ack => addr_of_2354_final_reg_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2354_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2354_request/$exit
      -- CP-element group 36: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2354_request/ack
      -- 
    ack_6845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2354_final_reg_ack_0, ack => convTransposeB_CP_6188_elements(36)); -- 
    -- CP-element group 37:  join  fork  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	85 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (24) 
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2354_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2354_complete/$exit
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2354_complete/ack
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_base_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_word_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_base_address_resized
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_base_addr_resize/$entry
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_base_addr_resize/$exit
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_base_addr_resize/base_resize_req
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_base_addr_resize/base_resize_ack
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_base_plus_offset/$entry
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_base_plus_offset/$exit
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_base_plus_offset/sum_rename_req
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_word_addrgen/$entry
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_word_addrgen/$exit
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_word_addrgen/root_register_req
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_word_addrgen/root_register_ack
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_Sample/word_access_start/$entry
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_Sample/word_access_start/word_0/$entry
      -- CP-element group 37: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_Sample/word_access_start/word_0/rr
      -- 
    ack_6850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2354_final_reg_ack_1, ack => convTransposeB_CP_6188_elements(37)); -- 
    rr_6883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(37), ack => ptr_deref_2358_load_0_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_Sample/word_access_start/$exit
      -- CP-element group 38: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_Sample/word_access_start/word_0/$exit
      -- CP-element group 38: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_Sample/word_access_start/word_0/ra
      -- 
    ra_6884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2358_load_0_ack_0, ack => convTransposeB_CP_6188_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	85 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	48 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_Update/word_access_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_Update/word_access_complete/word_0/$exit
      -- CP-element group 39: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_Update/word_access_complete/word_0/ca
      -- CP-element group 39: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_Update/ptr_deref_2358_Merge/$entry
      -- CP-element group 39: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_Update/ptr_deref_2358_Merge/$exit
      -- CP-element group 39: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_Update/ptr_deref_2358_Merge/merge_req
      -- CP-element group 39: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_Update/ptr_deref_2358_Merge/merge_ack
      -- 
    ca_6895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2358_load_0_ack_1, ack => convTransposeB_CP_6188_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	85 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2363_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2363_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2363_Sample/ra
      -- 
    ra_6909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2363_inst_ack_0, ack => convTransposeB_CP_6188_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	85 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2363_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2363_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2363_Update/ca
      -- CP-element group 41: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2377_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2377_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2377_Sample/rr
      -- 
    ca_6914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2363_inst_ack_1, ack => convTransposeB_CP_6188_elements(41)); -- 
    rr_6922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(41), ack => type_cast_2377_inst_req_0); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2377_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2377_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2377_Sample/ra
      -- 
    ra_6923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2377_inst_ack_0, ack => convTransposeB_CP_6188_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	85 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (16) 
      -- CP-element group 43: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_index_scale_1/$entry
      -- CP-element group 43: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2377_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2377_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2377_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_index_resized_1
      -- CP-element group 43: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_index_scaled_1
      -- CP-element group 43: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_index_computed_1
      -- CP-element group 43: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_index_resize_1/$entry
      -- CP-element group 43: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_index_resize_1/$exit
      -- CP-element group 43: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_index_resize_1/index_resize_req
      -- CP-element group 43: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_index_resize_1/index_resize_ack
      -- CP-element group 43: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_index_scale_1/$exit
      -- CP-element group 43: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_index_scale_1/scale_rename_req
      -- CP-element group 43: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_index_scale_1/scale_rename_ack
      -- CP-element group 43: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_final_index_sum_regn_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_final_index_sum_regn_Sample/req
      -- 
    ca_6928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2377_inst_ack_1, ack => convTransposeB_CP_6188_elements(43)); -- 
    req_6953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(43), ack => array_obj_ref_2383_index_offset_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	53 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_final_index_sum_regn_sample_complete
      -- CP-element group 44: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_final_index_sum_regn_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_final_index_sum_regn_Sample/ack
      -- 
    ack_6954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2383_index_offset_ack_0, ack => convTransposeB_CP_6188_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	85 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (11) 
      -- CP-element group 45: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2384_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_root_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_offset_calculated
      -- CP-element group 45: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_final_index_sum_regn_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_final_index_sum_regn_Update/ack
      -- CP-element group 45: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_base_plus_offset/$entry
      -- CP-element group 45: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_base_plus_offset/$exit
      -- CP-element group 45: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_base_plus_offset/sum_rename_req
      -- CP-element group 45: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_base_plus_offset/sum_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2384_request/$entry
      -- CP-element group 45: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2384_request/req
      -- 
    ack_6959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2383_index_offset_ack_1, ack => convTransposeB_CP_6188_elements(45)); -- 
    req_6968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(45), ack => addr_of_2384_final_reg_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2384_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2384_request/$exit
      -- CP-element group 46: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2384_request/ack
      -- 
    ack_6969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2384_final_reg_ack_0, ack => convTransposeB_CP_6188_elements(46)); -- 
    -- CP-element group 47:  fork  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	85 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (19) 
      -- CP-element group 47: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2384_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2384_complete/$exit
      -- CP-element group 47: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2384_complete/ack
      -- CP-element group 47: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_base_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_word_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_root_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_base_address_resized
      -- CP-element group 47: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_base_addr_resize/$entry
      -- CP-element group 47: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_base_addr_resize/$exit
      -- CP-element group 47: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_base_addr_resize/base_resize_req
      -- CP-element group 47: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_base_addr_resize/base_resize_ack
      -- CP-element group 47: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_base_plus_offset/$entry
      -- CP-element group 47: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_base_plus_offset/$exit
      -- CP-element group 47: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_base_plus_offset/sum_rename_req
      -- CP-element group 47: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_base_plus_offset/sum_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_word_addrgen/$entry
      -- CP-element group 47: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_word_addrgen/$exit
      -- CP-element group 47: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_word_addrgen/root_register_req
      -- CP-element group 47: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_word_addrgen/root_register_ack
      -- 
    ack_6974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2384_final_reg_ack_1, ack => convTransposeB_CP_6188_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: 	39 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (9) 
      -- CP-element group 48: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_Sample/ptr_deref_2387_Split/$entry
      -- CP-element group 48: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_Sample/ptr_deref_2387_Split/$exit
      -- CP-element group 48: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_Sample/ptr_deref_2387_Split/split_req
      -- CP-element group 48: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_Sample/ptr_deref_2387_Split/split_ack
      -- CP-element group 48: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_Sample/word_access_start/$entry
      -- CP-element group 48: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_Sample/word_access_start/word_0/$entry
      -- CP-element group 48: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_Sample/word_access_start/word_0/rr
      -- 
    rr_7012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(48), ack => ptr_deref_2387_store_0_req_0); -- 
    convTransposeB_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_6188_elements(47) & convTransposeB_CP_6188_elements(39);
      gj_convTransposeB_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_6188_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_Sample/word_access_start/$exit
      -- CP-element group 49: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_Sample/word_access_start/word_0/$exit
      -- CP-element group 49: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_Sample/word_access_start/word_0/ra
      -- 
    ra_7013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2387_store_0_ack_0, ack => convTransposeB_CP_6188_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	85 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_Update/word_access_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_Update/word_access_complete/word_0/$exit
      -- CP-element group 50: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_Update/word_access_complete/word_0/ca
      -- 
    ca_7024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2387_store_0_ack_1, ack => convTransposeB_CP_6188_elements(50)); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	85 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2393_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2393_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2393_Sample/ra
      -- 
    ra_7033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2393_inst_ack_0, ack => convTransposeB_CP_6188_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	85 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2393_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2393_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2393_Update/ca
      -- 
    ca_7038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2393_inst_ack_1, ack => convTransposeB_CP_6188_elements(52)); -- 
    -- CP-element group 53:  branch  join  transition  place  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	34 
    -- CP-element group 53: 	44 
    -- CP-element group 53: 	52 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (10) 
      -- CP-element group 53: 	 branch_block_stmt_2080/R_cmp_2409_place
      -- CP-element group 53: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407__exit__
      -- CP-element group 53: 	 branch_block_stmt_2080/if_stmt_2408__entry__
      -- CP-element group 53: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/$exit
      -- CP-element group 53: 	 branch_block_stmt_2080/if_stmt_2408_dead_link/$entry
      -- CP-element group 53: 	 branch_block_stmt_2080/if_stmt_2408_eval_test/$entry
      -- CP-element group 53: 	 branch_block_stmt_2080/if_stmt_2408_eval_test/$exit
      -- CP-element group 53: 	 branch_block_stmt_2080/if_stmt_2408_eval_test/branch_req
      -- CP-element group 53: 	 branch_block_stmt_2080/if_stmt_2408_if_link/$entry
      -- CP-element group 53: 	 branch_block_stmt_2080/if_stmt_2408_else_link/$entry
      -- 
    branch_req_7046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(53), ack => if_stmt_2408_branch_req_0); -- 
    convTransposeB_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_6188_elements(34) & convTransposeB_CP_6188_elements(44) & convTransposeB_CP_6188_elements(52) & convTransposeB_CP_6188_elements(50);
      gj_convTransposeB_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_6188_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	80 
    -- CP-element group 54: 	81 
    -- CP-element group 54:  members (24) 
      -- CP-element group 54: 	 branch_block_stmt_2080/whilex_xbody_ifx_xthen
      -- CP-element group 54: 	 branch_block_stmt_2080/merge_stmt_2414__exit__
      -- CP-element group 54: 	 branch_block_stmt_2080/assign_stmt_2420__entry__
      -- CP-element group 54: 	 branch_block_stmt_2080/assign_stmt_2420__exit__
      -- CP-element group 54: 	 branch_block_stmt_2080/ifx_xthen_whilex_xbody
      -- CP-element group 54: 	 branch_block_stmt_2080/if_stmt_2408_if_link/$exit
      -- CP-element group 54: 	 branch_block_stmt_2080/if_stmt_2408_if_link/if_choice_transition
      -- CP-element group 54: 	 branch_block_stmt_2080/assign_stmt_2420/$entry
      -- CP-element group 54: 	 branch_block_stmt_2080/assign_stmt_2420/$exit
      -- CP-element group 54: 	 branch_block_stmt_2080/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_2080/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2306/$entry
      -- CP-element group 54: 	 branch_block_stmt_2080/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2306/phi_stmt_2306_sources/$entry
      -- CP-element group 54: 	 branch_block_stmt_2080/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2306/phi_stmt_2306_sources/type_cast_2309/$entry
      -- CP-element group 54: 	 branch_block_stmt_2080/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2306/phi_stmt_2306_sources/type_cast_2309/SplitProtocol/$entry
      -- CP-element group 54: 	 branch_block_stmt_2080/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2306/phi_stmt_2306_sources/type_cast_2309/SplitProtocol/Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_2080/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2306/phi_stmt_2306_sources/type_cast_2309/SplitProtocol/Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_2080/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2306/phi_stmt_2306_sources/type_cast_2309/SplitProtocol/Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_2080/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2306/phi_stmt_2306_sources/type_cast_2309/SplitProtocol/Update/cr
      -- CP-element group 54: 	 branch_block_stmt_2080/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_2080/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 54: 	 branch_block_stmt_2080/merge_stmt_2414_PhiReqMerge
      -- CP-element group 54: 	 branch_block_stmt_2080/merge_stmt_2414_PhiAck/$entry
      -- CP-element group 54: 	 branch_block_stmt_2080/merge_stmt_2414_PhiAck/$exit
      -- CP-element group 54: 	 branch_block_stmt_2080/merge_stmt_2414_PhiAck/dummy
      -- 
    if_choice_transition_7051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2408_branch_ack_1, ack => convTransposeB_CP_6188_elements(54)); -- 
    rr_7235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(54), ack => type_cast_2309_inst_req_0); -- 
    cr_7240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(54), ack => type_cast_2309_inst_req_1); -- 
    -- CP-element group 55:  fork  transition  place  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	59 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (21) 
      -- CP-element group 55: 	 branch_block_stmt_2080/whilex_xbody_ifx_xelse
      -- CP-element group 55: 	 branch_block_stmt_2080/merge_stmt_2422__exit__
      -- CP-element group 55: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472__entry__
      -- CP-element group 55: 	 branch_block_stmt_2080/if_stmt_2408_else_link/$exit
      -- CP-element group 55: 	 branch_block_stmt_2080/if_stmt_2408_else_link/else_choice_transition
      -- CP-element group 55: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/$entry
      -- CP-element group 55: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2432_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2432_update_start_
      -- CP-element group 55: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2432_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2432_Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2432_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2432_Update/cr
      -- CP-element group 55: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2466_update_start_
      -- CP-element group 55: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2466_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2466_Update/cr
      -- CP-element group 55: 	 branch_block_stmt_2080/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 55: 	 branch_block_stmt_2080/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 55: 	 branch_block_stmt_2080/merge_stmt_2422_PhiReqMerge
      -- CP-element group 55: 	 branch_block_stmt_2080/merge_stmt_2422_PhiAck/$entry
      -- CP-element group 55: 	 branch_block_stmt_2080/merge_stmt_2422_PhiAck/$exit
      -- CP-element group 55: 	 branch_block_stmt_2080/merge_stmt_2422_PhiAck/dummy
      -- 
    else_choice_transition_7055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2408_branch_ack_0, ack => convTransposeB_CP_6188_elements(55)); -- 
    rr_7071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(55), ack => type_cast_2432_inst_req_0); -- 
    cr_7076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(55), ack => type_cast_2432_inst_req_1); -- 
    cr_7090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(55), ack => type_cast_2466_inst_req_1); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2432_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2432_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2432_Sample/ra
      -- 
    ra_7072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2432_inst_ack_0, ack => convTransposeB_CP_6188_elements(56)); -- 
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2432_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2432_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2432_Update/ca
      -- CP-element group 57: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2466_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2466_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2466_Sample/rr
      -- 
    ca_7077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2432_inst_ack_1, ack => convTransposeB_CP_6188_elements(57)); -- 
    rr_7085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(57), ack => type_cast_2466_inst_req_0); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2466_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2466_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2466_Sample/ra
      -- 
    ra_7086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2466_inst_ack_0, ack => convTransposeB_CP_6188_elements(58)); -- 
    -- CP-element group 59:  branch  transition  place  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	55 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (13) 
      -- CP-element group 59: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472__exit__
      -- CP-element group 59: 	 branch_block_stmt_2080/if_stmt_2473__entry__
      -- CP-element group 59: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/$exit
      -- CP-element group 59: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2466_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2466_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_2080/assign_stmt_2428_to_assign_stmt_2472/type_cast_2466_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_2080/if_stmt_2473_dead_link/$entry
      -- CP-element group 59: 	 branch_block_stmt_2080/if_stmt_2473_eval_test/$entry
      -- CP-element group 59: 	 branch_block_stmt_2080/if_stmt_2473_eval_test/$exit
      -- CP-element group 59: 	 branch_block_stmt_2080/if_stmt_2473_eval_test/branch_req
      -- CP-element group 59: 	 branch_block_stmt_2080/R_cmp100_2474_place
      -- CP-element group 59: 	 branch_block_stmt_2080/if_stmt_2473_if_link/$entry
      -- CP-element group 59: 	 branch_block_stmt_2080/if_stmt_2473_else_link/$entry
      -- 
    ca_7091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2466_inst_ack_1, ack => convTransposeB_CP_6188_elements(59)); -- 
    branch_req_7099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(59), ack => if_stmt_2473_branch_req_0); -- 
    -- CP-element group 60:  merge  transition  place  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (15) 
      -- CP-element group 60: 	 branch_block_stmt_2080/merge_stmt_2479__exit__
      -- CP-element group 60: 	 branch_block_stmt_2080/assign_stmt_2483__entry__
      -- CP-element group 60: 	 branch_block_stmt_2080/if_stmt_2473_if_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_2080/if_stmt_2473_if_link/if_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_2080/ifx_xelse_whilex_xend
      -- CP-element group 60: 	 branch_block_stmt_2080/assign_stmt_2483/$entry
      -- CP-element group 60: 	 branch_block_stmt_2080/assign_stmt_2483/WPIPE_Block1_done_2481_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2080/assign_stmt_2483/WPIPE_Block1_done_2481_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_2080/assign_stmt_2483/WPIPE_Block1_done_2481_Sample/req
      -- CP-element group 60: 	 branch_block_stmt_2080/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_2080/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_2080/merge_stmt_2479_PhiReqMerge
      -- CP-element group 60: 	 branch_block_stmt_2080/merge_stmt_2479_PhiAck/$entry
      -- CP-element group 60: 	 branch_block_stmt_2080/merge_stmt_2479_PhiAck/$exit
      -- CP-element group 60: 	 branch_block_stmt_2080/merge_stmt_2479_PhiAck/dummy
      -- 
    if_choice_transition_7104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2473_branch_ack_1, ack => convTransposeB_CP_6188_elements(60)); -- 
    req_7121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(60), ack => WPIPE_Block1_done_2481_inst_req_0); -- 
    -- CP-element group 61:  fork  transition  place  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	72 
    -- CP-element group 61: 	73 
    -- CP-element group 61: 	70 
    -- CP-element group 61: 	69 
    -- CP-element group 61:  members (20) 
      -- CP-element group 61: 	 branch_block_stmt_2080/if_stmt_2473_else_link/$exit
      -- CP-element group 61: 	 branch_block_stmt_2080/if_stmt_2473_else_link/else_choice_transition
      -- CP-element group 61: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 61: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/$entry
      -- CP-element group 61: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2245/$entry
      -- CP-element group 61: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2245/SplitProtocol/$entry
      -- CP-element group 61: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2245/SplitProtocol/Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2245/SplitProtocol/Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2245/SplitProtocol/Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2245/SplitProtocol/Update/cr
      -- CP-element group 61: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/$entry
      -- CP-element group 61: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/phi_stmt_2246_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/phi_stmt_2246_sources/type_cast_2252/$entry
      -- CP-element group 61: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/phi_stmt_2246_sources/type_cast_2252/SplitProtocol/$entry
      -- CP-element group 61: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/phi_stmt_2246_sources/type_cast_2252/SplitProtocol/Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/phi_stmt_2246_sources/type_cast_2252/SplitProtocol/Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/phi_stmt_2246_sources/type_cast_2252/SplitProtocol/Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/phi_stmt_2246_sources/type_cast_2252/SplitProtocol/Update/cr
      -- 
    else_choice_transition_7108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2473_branch_ack_0, ack => convTransposeB_CP_6188_elements(61)); -- 
    rr_7180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(61), ack => type_cast_2245_inst_req_0); -- 
    cr_7185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(61), ack => type_cast_2245_inst_req_1); -- 
    rr_7203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(61), ack => type_cast_2252_inst_req_0); -- 
    cr_7208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(61), ack => type_cast_2252_inst_req_1); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_2080/assign_stmt_2483/WPIPE_Block1_done_2481_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_2080/assign_stmt_2483/WPIPE_Block1_done_2481_update_start_
      -- CP-element group 62: 	 branch_block_stmt_2080/assign_stmt_2483/WPIPE_Block1_done_2481_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_2080/assign_stmt_2483/WPIPE_Block1_done_2481_Sample/ack
      -- CP-element group 62: 	 branch_block_stmt_2080/assign_stmt_2483/WPIPE_Block1_done_2481_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_2080/assign_stmt_2483/WPIPE_Block1_done_2481_Update/req
      -- 
    ack_7122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2481_inst_ack_0, ack => convTransposeB_CP_6188_elements(62)); -- 
    req_7126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(62), ack => WPIPE_Block1_done_2481_inst_req_1); -- 
    -- CP-element group 63:  transition  place  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (16) 
      -- CP-element group 63: 	 $exit
      -- CP-element group 63: 	 branch_block_stmt_2080/$exit
      -- CP-element group 63: 	 branch_block_stmt_2080/branch_block_stmt_2080__exit__
      -- CP-element group 63: 	 branch_block_stmt_2080/assign_stmt_2483__exit__
      -- CP-element group 63: 	 branch_block_stmt_2080/return__
      -- CP-element group 63: 	 branch_block_stmt_2080/merge_stmt_2485__exit__
      -- CP-element group 63: 	 branch_block_stmt_2080/assign_stmt_2483/$exit
      -- CP-element group 63: 	 branch_block_stmt_2080/assign_stmt_2483/WPIPE_Block1_done_2481_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_2080/assign_stmt_2483/WPIPE_Block1_done_2481_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_2080/assign_stmt_2483/WPIPE_Block1_done_2481_Update/ack
      -- CP-element group 63: 	 branch_block_stmt_2080/return___PhiReq/$entry
      -- CP-element group 63: 	 branch_block_stmt_2080/return___PhiReq/$exit
      -- CP-element group 63: 	 branch_block_stmt_2080/merge_stmt_2485_PhiReqMerge
      -- CP-element group 63: 	 branch_block_stmt_2080/merge_stmt_2485_PhiAck/$entry
      -- CP-element group 63: 	 branch_block_stmt_2080/merge_stmt_2485_PhiAck/$exit
      -- CP-element group 63: 	 branch_block_stmt_2080/merge_stmt_2485_PhiAck/dummy
      -- 
    ack_7127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2481_inst_ack_1, ack => convTransposeB_CP_6188_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	29 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/SplitProtocol/Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/SplitProtocol/Sample/ra
      -- 
    ra_7147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2243_inst_ack_0, ack => convTransposeB_CP_6188_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	29 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/SplitProtocol/Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/SplitProtocol/Update/ca
      -- 
    ca_7152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2243_inst_ack_1, ack => convTransposeB_CP_6188_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (5) 
      -- CP-element group 66: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/$exit
      -- CP-element group 66: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/$exit
      -- CP-element group 66: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/$exit
      -- CP-element group 66: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/SplitProtocol/$exit
      -- CP-element group 66: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_req
      -- 
    phi_stmt_2240_req_7153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2240_req_7153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(66), ack => phi_stmt_2240_req_0); -- 
    convTransposeB_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_6188_elements(65) & convTransposeB_CP_6188_elements(64);
      gj_convTransposeB_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_6188_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  transition  output  delay-element  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	29 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/$exit
      -- CP-element group 67: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/phi_stmt_2246_sources/$exit
      -- CP-element group 67: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/phi_stmt_2246_sources/type_cast_2250_konst_delay_trans
      -- CP-element group 67: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/phi_stmt_2246_req
      -- 
    phi_stmt_2246_req_7161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2246_req_7161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(67), ack => phi_stmt_2246_req_0); -- 
    -- Element group convTransposeB_CP_6188_elements(67) is a control-delay.
    cp_element_67_delay: control_delay_element  generic map(name => " 67_delay", delay_value => 1)  port map(req => convTransposeB_CP_6188_elements(29), ack => convTransposeB_CP_6188_elements(67), clk => clk, reset =>reset);
    -- CP-element group 68:  join  transition  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	76 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_2080/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_6188_elements(66) & convTransposeB_CP_6188_elements(67);
      gj_convTransposeB_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_6188_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	61 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2245/SplitProtocol/Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2245/SplitProtocol/Sample/ra
      -- 
    ra_7181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2245_inst_ack_0, ack => convTransposeB_CP_6188_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	61 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2245/SplitProtocol/Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2245/SplitProtocol/Update/ca
      -- 
    ca_7186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2245_inst_ack_1, ack => convTransposeB_CP_6188_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	75 
    -- CP-element group 71:  members (5) 
      -- CP-element group 71: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/$exit
      -- CP-element group 71: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/$exit
      -- CP-element group 71: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2245/$exit
      -- CP-element group 71: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2245/SplitProtocol/$exit
      -- CP-element group 71: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2240/phi_stmt_2240_req
      -- 
    phi_stmt_2240_req_7187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2240_req_7187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(71), ack => phi_stmt_2240_req_1); -- 
    convTransposeB_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_6188_elements(70) & convTransposeB_CP_6188_elements(69);
      gj_convTransposeB_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_6188_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	61 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/phi_stmt_2246_sources/type_cast_2252/SplitProtocol/Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/phi_stmt_2246_sources/type_cast_2252/SplitProtocol/Sample/ra
      -- 
    ra_7204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2252_inst_ack_0, ack => convTransposeB_CP_6188_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	61 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/phi_stmt_2246_sources/type_cast_2252/SplitProtocol/Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/phi_stmt_2246_sources/type_cast_2252/SplitProtocol/Update/ca
      -- 
    ca_7209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2252_inst_ack_1, ack => convTransposeB_CP_6188_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/$exit
      -- CP-element group 74: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/phi_stmt_2246_sources/$exit
      -- CP-element group 74: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/phi_stmt_2246_sources/type_cast_2252/$exit
      -- CP-element group 74: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/phi_stmt_2246_sources/type_cast_2252/SplitProtocol/$exit
      -- CP-element group 74: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2246/phi_stmt_2246_req
      -- 
    phi_stmt_2246_req_7210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2246_req_7210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(74), ack => phi_stmt_2246_req_1); -- 
    convTransposeB_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_6188_elements(72) & convTransposeB_CP_6188_elements(73);
      gj_convTransposeB_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_6188_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: 	71 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_2080/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_6188_elements(74) & convTransposeB_CP_6188_elements(71);
      gj_convTransposeB_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_6188_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  merge  fork  transition  place  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: 	68 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_2080/merge_stmt_2239_PhiReqMerge
      -- CP-element group 76: 	 branch_block_stmt_2080/merge_stmt_2239_PhiAck/$entry
      -- 
    convTransposeB_CP_6188_elements(76) <= OrReduce(convTransposeB_CP_6188_elements(75) & convTransposeB_CP_6188_elements(68));
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_2080/merge_stmt_2239_PhiAck/phi_stmt_2240_ack
      -- 
    phi_stmt_2240_ack_7215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2240_ack_0, ack => convTransposeB_CP_6188_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_2080/merge_stmt_2239_PhiAck/phi_stmt_2246_ack
      -- 
    phi_stmt_2246_ack_7216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2246_ack_0, ack => convTransposeB_CP_6188_elements(78)); -- 
    -- CP-element group 79:  join  transition  place  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	83 
    -- CP-element group 79:  members (10) 
      -- CP-element group 79: 	 branch_block_stmt_2080/merge_stmt_2239__exit__
      -- CP-element group 79: 	 branch_block_stmt_2080/assign_stmt_2258_to_assign_stmt_2303__entry__
      -- CP-element group 79: 	 branch_block_stmt_2080/assign_stmt_2258_to_assign_stmt_2303__exit__
      -- CP-element group 79: 	 branch_block_stmt_2080/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 79: 	 branch_block_stmt_2080/assign_stmt_2258_to_assign_stmt_2303/$entry
      -- CP-element group 79: 	 branch_block_stmt_2080/assign_stmt_2258_to_assign_stmt_2303/$exit
      -- CP-element group 79: 	 branch_block_stmt_2080/merge_stmt_2239_PhiAck/$exit
      -- CP-element group 79: 	 branch_block_stmt_2080/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 79: 	 branch_block_stmt_2080/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2306/$entry
      -- CP-element group 79: 	 branch_block_stmt_2080/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2306/phi_stmt_2306_sources/$entry
      -- 
    convTransposeB_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_6188_elements(77) & convTransposeB_CP_6188_elements(78);
      gj_convTransposeB_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_6188_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	54 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_2080/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2306/phi_stmt_2306_sources/type_cast_2309/SplitProtocol/Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_2080/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2306/phi_stmt_2306_sources/type_cast_2309/SplitProtocol/Sample/ra
      -- 
    ra_7236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2309_inst_ack_0, ack => convTransposeB_CP_6188_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	54 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_2080/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2306/phi_stmt_2306_sources/type_cast_2309/SplitProtocol/Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_2080/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2306/phi_stmt_2306_sources/type_cast_2309/SplitProtocol/Update/ca
      -- 
    ca_7241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2309_inst_ack_1, ack => convTransposeB_CP_6188_elements(81)); -- 
    -- CP-element group 82:  join  transition  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_2080/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 82: 	 branch_block_stmt_2080/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2306/$exit
      -- CP-element group 82: 	 branch_block_stmt_2080/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2306/phi_stmt_2306_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_2080/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2306/phi_stmt_2306_sources/type_cast_2309/$exit
      -- CP-element group 82: 	 branch_block_stmt_2080/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2306/phi_stmt_2306_sources/type_cast_2309/SplitProtocol/$exit
      -- CP-element group 82: 	 branch_block_stmt_2080/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2306/phi_stmt_2306_req
      -- 
    phi_stmt_2306_req_7242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2306_req_7242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(82), ack => phi_stmt_2306_req_0); -- 
    convTransposeB_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_6188_elements(80) & convTransposeB_CP_6188_elements(81);
      gj_convTransposeB_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_6188_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  transition  output  delay-element  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	79 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (5) 
      -- CP-element group 83: 	 branch_block_stmt_2080/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 83: 	 branch_block_stmt_2080/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2306/$exit
      -- CP-element group 83: 	 branch_block_stmt_2080/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2306/phi_stmt_2306_sources/$exit
      -- CP-element group 83: 	 branch_block_stmt_2080/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2306/phi_stmt_2306_sources/type_cast_2312_konst_delay_trans
      -- CP-element group 83: 	 branch_block_stmt_2080/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2306/phi_stmt_2306_req
      -- 
    phi_stmt_2306_req_7253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2306_req_7253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(83), ack => phi_stmt_2306_req_1); -- 
    -- Element group convTransposeB_CP_6188_elements(83) is a control-delay.
    cp_element_83_delay: control_delay_element  generic map(name => " 83_delay", delay_value => 1)  port map(req => convTransposeB_CP_6188_elements(79), ack => convTransposeB_CP_6188_elements(83), clk => clk, reset =>reset);
    -- CP-element group 84:  merge  transition  place  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_2080/merge_stmt_2305_PhiReqMerge
      -- CP-element group 84: 	 branch_block_stmt_2080/merge_stmt_2305_PhiAck/$entry
      -- 
    convTransposeB_CP_6188_elements(84) <= OrReduce(convTransposeB_CP_6188_elements(82) & convTransposeB_CP_6188_elements(83));
    -- CP-element group 85:  fork  transition  place  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	30 
    -- CP-element group 85: 	31 
    -- CP-element group 85: 	35 
    -- CP-element group 85: 	45 
    -- CP-element group 85: 	37 
    -- CP-element group 85: 	51 
    -- CP-element group 85: 	52 
    -- CP-element group 85: 	47 
    -- CP-element group 85: 	40 
    -- CP-element group 85: 	41 
    -- CP-element group 85: 	50 
    -- CP-element group 85: 	39 
    -- CP-element group 85: 	43 
    -- CP-element group 85: 	33 
    -- CP-element group 85:  members (51) 
      -- CP-element group 85: 	 branch_block_stmt_2080/merge_stmt_2305__exit__
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407__entry__
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/$entry
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2333_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2333_update_start_
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2333_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2333_Sample/rr
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2333_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2333_Update/cr
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2347_update_start_
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2347_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2347_Update/cr
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2354_update_start_
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_final_index_sum_regn_update_start
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_final_index_sum_regn_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2353_final_index_sum_regn_Update/req
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2354_complete/$entry
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2354_complete/req
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_update_start_
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_Update/word_access_complete/$entry
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_Update/word_access_complete/word_0/$entry
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2358_Update/word_access_complete/word_0/cr
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2363_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2363_update_start_
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2363_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2363_Sample/rr
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2363_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2363_Update/cr
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2377_update_start_
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2377_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2377_Update/cr
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2384_update_start_
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_final_index_sum_regn_update_start
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_final_index_sum_regn_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/array_obj_ref_2383_final_index_sum_regn_Update/req
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2384_complete/$entry
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/addr_of_2384_complete/req
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_update_start_
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_Update/word_access_complete/$entry
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_Update/word_access_complete/word_0/$entry
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/ptr_deref_2387_Update/word_access_complete/word_0/cr
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2393_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2393_update_start_
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2393_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2393_Sample/rr
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2393_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_2080/assign_stmt_2319_to_assign_stmt_2407/type_cast_2393_Update/cr
      -- CP-element group 85: 	 branch_block_stmt_2080/merge_stmt_2305_PhiAck/$exit
      -- CP-element group 85: 	 branch_block_stmt_2080/merge_stmt_2305_PhiAck/phi_stmt_2306_ack
      -- 
    phi_stmt_2306_ack_7258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2306_ack_0, ack => convTransposeB_CP_6188_elements(85)); -- 
    rr_6784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(85), ack => type_cast_2333_inst_req_0); -- 
    cr_6789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(85), ack => type_cast_2333_inst_req_1); -- 
    cr_6803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(85), ack => type_cast_2347_inst_req_1); -- 
    req_6834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(85), ack => array_obj_ref_2353_index_offset_req_1); -- 
    req_6849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(85), ack => addr_of_2354_final_reg_req_1); -- 
    cr_6894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(85), ack => ptr_deref_2358_load_0_req_1); -- 
    rr_6908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(85), ack => type_cast_2363_inst_req_0); -- 
    cr_6913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(85), ack => type_cast_2363_inst_req_1); -- 
    cr_6927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(85), ack => type_cast_2377_inst_req_1); -- 
    req_6958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(85), ack => array_obj_ref_2383_index_offset_req_1); -- 
    req_6973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(85), ack => addr_of_2384_final_reg_req_1); -- 
    cr_7023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(85), ack => ptr_deref_2387_store_0_req_1); -- 
    rr_7032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(85), ack => type_cast_2393_inst_req_0); -- 
    cr_7037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_6188_elements(85), ack => type_cast_2393_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2341_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2371_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_2138_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_2138_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom68_2382_resized : std_logic_vector(13 downto 0);
    signal R_idxprom68_2382_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2352_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2352_scaled : std_logic_vector(13 downto 0);
    signal add20_2324 : std_logic_vector(15 downto 0);
    signal add60_2329 : std_logic_vector(15 downto 0);
    signal add73_2400 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2353_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2353_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2353_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2353_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2353_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2353_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2383_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2383_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2383_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2383_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2383_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2383_root_address : std_logic_vector(13 downto 0);
    signal arrayidx69_2385 : std_logic_vector(31 downto 0);
    signal arrayidx_2355 : std_logic_vector(31 downto 0);
    signal call_2083 : std_logic_vector(15 downto 0);
    signal cmp100_2472 : std_logic_vector(0 downto 0);
    signal cmp86_2438 : std_logic_vector(0 downto 0);
    signal cmp_2407 : std_logic_vector(0 downto 0);
    signal conv63_2334 : std_logic_vector(31 downto 0);
    signal conv66_2364 : std_logic_vector(31 downto 0);
    signal conv72_2394 : std_logic_vector(31 downto 0);
    signal conv75_2189 : std_logic_vector(31 downto 0);
    signal conv83_2433 : std_logic_vector(31 downto 0);
    signal conv85_2193 : std_logic_vector(31 downto 0);
    signal conv96_2467 : std_logic_vector(31 downto 0);
    signal conv98_2209 : std_logic_vector(31 downto 0);
    signal div93_2450 : std_logic_vector(15 downto 0);
    signal div99_2215 : std_logic_vector(31 downto 0);
    signal div_2102 : std_logic_vector(15 downto 0);
    signal iNsTr_10_2201 : std_logic_vector(31 downto 0);
    signal iNsTr_2_2092 : std_logic_vector(31 downto 0);
    signal iNsTr_3_2110 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2120 : std_logic_vector(31 downto 0);
    signal iNsTr_5_2132 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2145 : std_logic_vector(31 downto 0);
    signal iNsTr_7_2157 : std_logic_vector(31 downto 0);
    signal iNsTr_8_2169 : std_logic_vector(31 downto 0);
    signal iNsTr_9_2181 : std_logic_vector(31 downto 0);
    signal idxprom68_2378 : std_logic_vector(63 downto 0);
    signal idxprom_2348 : std_logic_vector(63 downto 0);
    signal inc90_2444 : std_logic_vector(15 downto 0);
    signal inc_2428 : std_logic_vector(15 downto 0);
    signal indvar_2306 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2420 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_2462 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2246 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2240 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2456 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2319 : std_logic_vector(15 downto 0);
    signal ptr_deref_2095_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2095_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2095_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2095_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2095_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2113_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2113_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2113_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2113_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2113_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2123_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2123_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2123_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2123_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2123_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2135_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2135_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2135_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2135_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2135_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2148_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2148_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2148_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2148_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2148_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2160_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2160_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2160_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2160_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2160_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2172_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2172_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2172_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2172_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2172_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2184_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2184_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2184_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2184_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2184_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2204_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2204_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2204_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2204_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2204_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2358_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2358_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2358_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2358_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2358_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2387_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2387_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2387_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2387_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2387_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2387_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr67_2373 : std_logic_vector(31 downto 0);
    signal shr_2343 : std_logic_vector(31 downto 0);
    signal tmp10_2288 : std_logic_vector(15 downto 0);
    signal tmp11_2114 : std_logic_vector(15 downto 0);
    signal tmp128_2258 : std_logic_vector(15 downto 0);
    signal tmp129_2263 : std_logic_vector(15 downto 0);
    signal tmp12_2293 : std_logic_vector(15 downto 0);
    signal tmp130_2268 : std_logic_vector(15 downto 0);
    signal tmp13_2298 : std_logic_vector(15 downto 0);
    signal tmp14_2303 : std_logic_vector(15 downto 0);
    signal tmp24_2124 : std_logic_vector(15 downto 0);
    signal tmp27_2136 : std_logic_vector(15 downto 0);
    signal tmp30_2139 : std_logic_vector(15 downto 0);
    signal tmp36_2149 : std_logic_vector(15 downto 0);
    signal tmp39_2161 : std_logic_vector(15 downto 0);
    signal tmp3_2221 : std_logic_vector(15 downto 0);
    signal tmp49_2173 : std_logic_vector(15 downto 0);
    signal tmp4_2226 : std_logic_vector(15 downto 0);
    signal tmp53_2185 : std_logic_vector(15 downto 0);
    signal tmp5_2273 : std_logic_vector(15 downto 0);
    signal tmp64_2359 : std_logic_vector(63 downto 0);
    signal tmp6_2278 : std_logic_vector(15 downto 0);
    signal tmp7_2232 : std_logic_vector(15 downto 0);
    signal tmp8_2237 : std_logic_vector(15 downto 0);
    signal tmp97_2205 : std_logic_vector(15 downto 0);
    signal tmp9_2283 : std_logic_vector(15 downto 0);
    signal tmp_2096 : std_logic_vector(15 downto 0);
    signal type_cast_2100_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2213_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2219_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2230_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2243_wire : std_logic_vector(15 downto 0);
    signal type_cast_2245_wire : std_logic_vector(15 downto 0);
    signal type_cast_2250_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2252_wire : std_logic_vector(15 downto 0);
    signal type_cast_2309_wire : std_logic_vector(15 downto 0);
    signal type_cast_2312_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2317_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2332_wire : std_logic_vector(31 downto 0);
    signal type_cast_2337_wire : std_logic_vector(31 downto 0);
    signal type_cast_2340_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2346_wire : std_logic_vector(63 downto 0);
    signal type_cast_2362_wire : std_logic_vector(31 downto 0);
    signal type_cast_2367_wire : std_logic_vector(31 downto 0);
    signal type_cast_2370_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2376_wire : std_logic_vector(63 downto 0);
    signal type_cast_2392_wire : std_logic_vector(31 downto 0);
    signal type_cast_2398_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2403_wire : std_logic_vector(31 downto 0);
    signal type_cast_2405_wire : std_logic_vector(31 downto 0);
    signal type_cast_2418_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2426_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2431_wire : std_logic_vector(31 downto 0);
    signal type_cast_2442_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2448_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2465_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_2138_word_address_0 <= "0";
    array_obj_ref_2353_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2353_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2353_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2353_resized_base_address <= "00000000000000";
    array_obj_ref_2383_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2383_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2383_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2383_resized_base_address <= "00000000000000";
    iNsTr_10_2201 <= "00000000000000000000000000000100";
    iNsTr_2_2092 <= "00000000000000000000000000000101";
    iNsTr_3_2110 <= "00000000000000000000000000000110";
    iNsTr_4_2120 <= "00000000000000000000000000000000";
    iNsTr_5_2132 <= "00000000000000000000000000000101";
    iNsTr_6_2145 <= "00000000000000000000000000000001";
    iNsTr_7_2157 <= "00000000000000000000000000000110";
    iNsTr_8_2169 <= "00000000000000000000000000000110";
    iNsTr_9_2181 <= "00000000000000000000000000000101";
    ptr_deref_2095_word_offset_0 <= "0000000";
    ptr_deref_2113_word_offset_0 <= "0000000";
    ptr_deref_2123_word_offset_0 <= "0";
    ptr_deref_2135_word_offset_0 <= "0000000";
    ptr_deref_2148_word_offset_0 <= "0";
    ptr_deref_2160_word_offset_0 <= "0000000";
    ptr_deref_2172_word_offset_0 <= "0000000";
    ptr_deref_2184_word_offset_0 <= "0000000";
    ptr_deref_2204_word_offset_0 <= "0000000";
    ptr_deref_2358_word_offset_0 <= "00000000000000";
    ptr_deref_2387_word_offset_0 <= "00000000000000";
    type_cast_2100_wire_constant <= "0000000000000001";
    type_cast_2213_wire_constant <= "00000000000000000000000000000001";
    type_cast_2219_wire_constant <= "1111111111111111";
    type_cast_2230_wire_constant <= "1111111111111111";
    type_cast_2250_wire_constant <= "0000000000000000";
    type_cast_2312_wire_constant <= "0000000000000000";
    type_cast_2317_wire_constant <= "0000000000000100";
    type_cast_2340_wire_constant <= "00000000000000000000000000000010";
    type_cast_2370_wire_constant <= "00000000000000000000000000000010";
    type_cast_2398_wire_constant <= "00000000000000000000000000000100";
    type_cast_2418_wire_constant <= "0000000000000001";
    type_cast_2426_wire_constant <= "0000000000000001";
    type_cast_2442_wire_constant <= "0000000000000001";
    type_cast_2448_wire_constant <= "0000000000000001";
    phi_stmt_2240: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2243_wire & type_cast_2245_wire;
      req <= phi_stmt_2240_req_0 & phi_stmt_2240_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2240",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2240_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2240,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2240
    phi_stmt_2246: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2250_wire_constant & type_cast_2252_wire;
      req <= phi_stmt_2246_req_0 & phi_stmt_2246_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2246",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2246_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2246,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2246
    phi_stmt_2306: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2309_wire & type_cast_2312_wire_constant;
      req <= phi_stmt_2306_req_0 & phi_stmt_2306_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2306",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2306_ack_0,
          idata => idata,
          odata => indvar_2306,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2306
    -- flow-through select operator MUX_2455_inst
    input_dim1x_x2_2456 <= div93_2450 when (cmp86_2438(0) /=  '0') else inc_2428;
    -- flow-through select operator MUX_2461_inst
    input_dim0x_x0_2462 <= inc90_2444 when (cmp86_2438(0) /=  '0') else input_dim0x_x2x_xph_2246;
    addr_of_2354_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2354_final_reg_req_0;
      addr_of_2354_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2354_final_reg_req_1;
      addr_of_2354_final_reg_ack_1<= rack(0);
      addr_of_2354_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2354_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2353_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_2355,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2384_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2384_final_reg_req_0;
      addr_of_2384_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2384_final_reg_req_1;
      addr_of_2384_final_reg_ack_1<= rack(0);
      addr_of_2384_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2384_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2383_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx69_2385,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2188_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2188_inst_req_0;
      type_cast_2188_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2188_inst_req_1;
      type_cast_2188_inst_ack_1<= rack(0);
      type_cast_2188_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2188_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp11_2114,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2189,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2192_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2192_inst_req_0;
      type_cast_2192_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2192_inst_req_1;
      type_cast_2192_inst_ack_1<= rack(0);
      type_cast_2192_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2192_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_2096,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_2193,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2208_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2208_inst_req_0;
      type_cast_2208_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2208_inst_req_1;
      type_cast_2208_inst_ack_1<= rack(0);
      type_cast_2208_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2208_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp97_2205,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_2209,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2243_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2243_inst_req_0;
      type_cast_2243_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2243_inst_req_1;
      type_cast_2243_inst_ack_1<= rack(0);
      type_cast_2243_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2243_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2102,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2243_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2245_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2245_inst_req_0;
      type_cast_2245_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2245_inst_req_1;
      type_cast_2245_inst_ack_1<= rack(0);
      type_cast_2245_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2245_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2456,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2245_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2252_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2252_inst_req_0;
      type_cast_2252_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2252_inst_req_1;
      type_cast_2252_inst_ack_1<= rack(0);
      type_cast_2252_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2252_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_2462,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2252_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2309_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2309_inst_req_0;
      type_cast_2309_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2309_inst_req_1;
      type_cast_2309_inst_ack_1<= rack(0);
      type_cast_2309_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2309_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2420,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2309_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2333_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2333_inst_req_0;
      type_cast_2333_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2333_inst_req_1;
      type_cast_2333_inst_ack_1<= rack(0);
      type_cast_2333_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2333_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2332_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_2334,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2337_inst
    process(conv63_2334) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv63_2334(31 downto 0);
      type_cast_2337_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2342_inst
    process(ASHR_i32_i32_2341_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2341_wire(31 downto 0);
      shr_2343 <= tmp_var; -- 
    end process;
    type_cast_2347_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2347_inst_req_0;
      type_cast_2347_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2347_inst_req_1;
      type_cast_2347_inst_ack_1<= rack(0);
      type_cast_2347_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2347_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2346_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2348,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2363_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2363_inst_req_0;
      type_cast_2363_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2363_inst_req_1;
      type_cast_2363_inst_ack_1<= rack(0);
      type_cast_2363_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2363_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2362_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_2364,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2367_inst
    process(conv66_2364) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv66_2364(31 downto 0);
      type_cast_2367_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2372_inst
    process(ASHR_i32_i32_2371_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2371_wire(31 downto 0);
      shr67_2373 <= tmp_var; -- 
    end process;
    type_cast_2377_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2377_inst_req_0;
      type_cast_2377_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2377_inst_req_1;
      type_cast_2377_inst_ack_1<= rack(0);
      type_cast_2377_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2377_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2376_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom68_2378,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2393_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2393_inst_req_0;
      type_cast_2393_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2393_inst_req_1;
      type_cast_2393_inst_ack_1<= rack(0);
      type_cast_2393_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2393_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2392_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv72_2394,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2403_inst
    process(add73_2400) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add73_2400(31 downto 0);
      type_cast_2403_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2405_inst
    process(conv75_2189) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv75_2189(31 downto 0);
      type_cast_2405_wire <= tmp_var; -- 
    end process;
    type_cast_2432_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2432_inst_req_0;
      type_cast_2432_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2432_inst_req_1;
      type_cast_2432_inst_ack_1<= rack(0);
      type_cast_2432_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2432_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2431_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_2433,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2466_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2466_inst_req_0;
      type_cast_2466_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2466_inst_req_1;
      type_cast_2466_inst_ack_1<= rack(0);
      type_cast_2466_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2466_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2465_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv96_2467,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_2138_gather_scatter
    process(LOAD_padding_2138_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_2138_data_0;
      ov(15 downto 0) := iv;
      tmp30_2139 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2353_index_1_rename
    process(R_idxprom_2352_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2352_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2352_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2353_index_1_resize
    process(idxprom_2348) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2348;
      ov := iv(13 downto 0);
      R_idxprom_2352_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2353_root_address_inst
    process(array_obj_ref_2353_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2353_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2353_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2383_index_1_rename
    process(R_idxprom68_2382_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom68_2382_resized;
      ov(13 downto 0) := iv;
      R_idxprom68_2382_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2383_index_1_resize
    process(idxprom68_2378) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom68_2378;
      ov := iv(13 downto 0);
      R_idxprom68_2382_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2383_root_address_inst
    process(array_obj_ref_2383_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2383_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2383_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2095_addr_0
    process(ptr_deref_2095_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2095_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2095_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2095_base_resize
    process(iNsTr_2_2092) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_2092;
      ov := iv(6 downto 0);
      ptr_deref_2095_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2095_gather_scatter
    process(ptr_deref_2095_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2095_data_0;
      ov(15 downto 0) := iv;
      tmp_2096 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2095_root_address_inst
    process(ptr_deref_2095_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2095_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2095_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2113_addr_0
    process(ptr_deref_2113_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2113_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2113_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2113_base_resize
    process(iNsTr_3_2110) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_2110;
      ov := iv(6 downto 0);
      ptr_deref_2113_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2113_gather_scatter
    process(ptr_deref_2113_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2113_data_0;
      ov(15 downto 0) := iv;
      tmp11_2114 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2113_root_address_inst
    process(ptr_deref_2113_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2113_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2113_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2123_addr_0
    process(ptr_deref_2123_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2123_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2123_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2123_base_resize
    process(iNsTr_4_2120) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_2120;
      ov := iv(0 downto 0);
      ptr_deref_2123_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2123_gather_scatter
    process(ptr_deref_2123_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2123_data_0;
      ov(15 downto 0) := iv;
      tmp24_2124 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2123_root_address_inst
    process(ptr_deref_2123_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2123_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2123_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2135_addr_0
    process(ptr_deref_2135_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2135_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2135_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2135_base_resize
    process(iNsTr_5_2132) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_2132;
      ov := iv(6 downto 0);
      ptr_deref_2135_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2135_gather_scatter
    process(ptr_deref_2135_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2135_data_0;
      ov(15 downto 0) := iv;
      tmp27_2136 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2135_root_address_inst
    process(ptr_deref_2135_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2135_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2135_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2148_addr_0
    process(ptr_deref_2148_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2148_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2148_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2148_base_resize
    process(iNsTr_6_2145) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_2145;
      ov := iv(0 downto 0);
      ptr_deref_2148_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2148_gather_scatter
    process(ptr_deref_2148_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2148_data_0;
      ov(15 downto 0) := iv;
      tmp36_2149 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2148_root_address_inst
    process(ptr_deref_2148_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2148_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2148_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2160_addr_0
    process(ptr_deref_2160_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2160_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2160_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2160_base_resize
    process(iNsTr_7_2157) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_2157;
      ov := iv(6 downto 0);
      ptr_deref_2160_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2160_gather_scatter
    process(ptr_deref_2160_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2160_data_0;
      ov(15 downto 0) := iv;
      tmp39_2161 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2160_root_address_inst
    process(ptr_deref_2160_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2160_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2160_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2172_addr_0
    process(ptr_deref_2172_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2172_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2172_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2172_base_resize
    process(iNsTr_8_2169) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_2169;
      ov := iv(6 downto 0);
      ptr_deref_2172_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2172_gather_scatter
    process(ptr_deref_2172_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2172_data_0;
      ov(15 downto 0) := iv;
      tmp49_2173 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2172_root_address_inst
    process(ptr_deref_2172_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2172_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2172_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2184_addr_0
    process(ptr_deref_2184_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2184_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2184_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2184_base_resize
    process(iNsTr_9_2181) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_2181;
      ov := iv(6 downto 0);
      ptr_deref_2184_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2184_gather_scatter
    process(ptr_deref_2184_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2184_data_0;
      ov(15 downto 0) := iv;
      tmp53_2185 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2184_root_address_inst
    process(ptr_deref_2184_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2184_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2184_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2204_addr_0
    process(ptr_deref_2204_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2204_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2204_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2204_base_resize
    process(iNsTr_10_2201) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_2201;
      ov := iv(6 downto 0);
      ptr_deref_2204_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2204_gather_scatter
    process(ptr_deref_2204_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2204_data_0;
      ov(15 downto 0) := iv;
      tmp97_2205 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2204_root_address_inst
    process(ptr_deref_2204_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2204_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2204_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2358_addr_0
    process(ptr_deref_2358_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2358_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2358_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2358_base_resize
    process(arrayidx_2355) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_2355;
      ov := iv(13 downto 0);
      ptr_deref_2358_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2358_gather_scatter
    process(ptr_deref_2358_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2358_data_0;
      ov(63 downto 0) := iv;
      tmp64_2359 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2358_root_address_inst
    process(ptr_deref_2358_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2358_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2358_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2387_addr_0
    process(ptr_deref_2387_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2387_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2387_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2387_base_resize
    process(arrayidx69_2385) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx69_2385;
      ov := iv(13 downto 0);
      ptr_deref_2387_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2387_gather_scatter
    process(tmp64_2359) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp64_2359;
      ov(63 downto 0) := iv;
      ptr_deref_2387_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2387_root_address_inst
    process(ptr_deref_2387_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2387_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2387_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2408_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2407;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2408_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2408_branch_req_0,
          ack0 => if_stmt_2408_branch_ack_0,
          ack1 => if_stmt_2408_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2473_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp100_2472;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2473_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2473_branch_req_0,
          ack0 => if_stmt_2473_branch_ack_0,
          ack1 => if_stmt_2473_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2220_inst
    process(tmp39_2161) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp39_2161, type_cast_2219_wire_constant, tmp_var);
      tmp3_2221 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2231_inst
    process(tmp27_2136) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp27_2136, type_cast_2230_wire_constant, tmp_var);
      tmp7_2232 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2262_inst
    process(input_dim1x_x1x_xph_2240, tmp128_2258) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2240, tmp128_2258, tmp_var);
      tmp129_2263 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2277_inst
    process(tmp4_2226, tmp5_2273) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp4_2226, tmp5_2273, tmp_var);
      tmp6_2278 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2287_inst
    process(tmp8_2237, tmp9_2283) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp8_2237, tmp9_2283, tmp_var);
      tmp10_2288 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2297_inst
    process(tmp6_2278, tmp12_2293) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp6_2278, tmp12_2293, tmp_var);
      tmp13_2298 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2323_inst
    process(tmp130_2268, input_dim2x_x1_2319) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp130_2268, input_dim2x_x1_2319, tmp_var);
      add20_2324 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2328_inst
    process(tmp14_2303, input_dim2x_x1_2319) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp14_2303, input_dim2x_x1_2319, tmp_var);
      add60_2329 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2419_inst
    process(indvar_2306) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2306, type_cast_2418_wire_constant, tmp_var);
      indvarx_xnext_2420 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2427_inst
    process(input_dim1x_x1x_xph_2240) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2240, type_cast_2426_wire_constant, tmp_var);
      inc_2428 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2443_inst
    process(input_dim0x_x2x_xph_2246) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim0x_x2x_xph_2246, type_cast_2442_wire_constant, tmp_var);
      inc90_2444 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2399_inst
    process(conv72_2394) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv72_2394, type_cast_2398_wire_constant, tmp_var);
      add73_2400 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2341_inst
    process(type_cast_2337_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2337_wire, type_cast_2340_wire_constant, tmp_var);
      ASHR_i32_i32_2341_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2371_inst
    process(type_cast_2367_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2367_wire, type_cast_2370_wire_constant, tmp_var);
      ASHR_i32_i32_2371_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2437_inst
    process(conv83_2433, conv85_2193) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv83_2433, conv85_2193, tmp_var);
      cmp86_2438 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2471_inst
    process(conv96_2467, div99_2215) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv96_2467, div99_2215, tmp_var);
      cmp100_2472 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2101_inst
    process(tmp_2096) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_2096, type_cast_2100_wire_constant, tmp_var);
      div_2102 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2449_inst
    process(tmp_2096) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_2096, type_cast_2448_wire_constant, tmp_var);
      div93_2450 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2214_inst
    process(conv98_2209) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv98_2209, type_cast_2213_wire_constant, tmp_var);
      div99_2215 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2257_inst
    process(tmp_2096, input_dim0x_x2x_xph_2246) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp_2096, input_dim0x_x2x_xph_2246, tmp_var);
      tmp128_2258 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2267_inst
    process(tmp11_2114, tmp129_2263) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp11_2114, tmp129_2263, tmp_var);
      tmp130_2268 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2272_inst
    process(tmp36_2149, input_dim1x_x1x_xph_2240) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp36_2149, input_dim1x_x1x_xph_2240, tmp_var);
      tmp5_2273 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2282_inst
    process(tmp24_2124, input_dim0x_x2x_xph_2246) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp24_2124, input_dim0x_x2x_xph_2246, tmp_var);
      tmp9_2283 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2292_inst
    process(tmp53_2185, tmp10_2288) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp53_2185, tmp10_2288, tmp_var);
      tmp12_2293 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2302_inst
    process(tmp49_2173, tmp13_2298) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp49_2173, tmp13_2298, tmp_var);
      tmp14_2303 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2318_inst
    process(indvar_2306) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2306, type_cast_2317_wire_constant, tmp_var);
      input_dim2x_x1_2319 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2406_inst
    process(type_cast_2403_wire, type_cast_2405_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2403_wire, type_cast_2405_wire, tmp_var);
      cmp_2407 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2225_inst
    process(tmp3_2221, tmp30_2139) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp3_2221, tmp30_2139, tmp_var);
      tmp4_2226 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2236_inst
    process(tmp7_2232, tmp30_2139) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp7_2232, tmp30_2139, tmp_var);
      tmp8_2237 <= tmp_var; --
    end process;
    -- shared split operator group (29) : array_obj_ref_2353_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2352_scaled;
      array_obj_ref_2353_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2353_index_offset_req_0;
      array_obj_ref_2353_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2353_index_offset_req_1;
      array_obj_ref_2353_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : array_obj_ref_2383_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom68_2382_scaled;
      array_obj_ref_2383_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2383_index_offset_req_0;
      array_obj_ref_2383_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2383_index_offset_req_1;
      array_obj_ref_2383_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- unary operator type_cast_2332_inst
    process(add20_2324) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add20_2324, tmp_var);
      type_cast_2332_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2346_inst
    process(shr_2343) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2343, tmp_var);
      type_cast_2346_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2362_inst
    process(add60_2329) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add60_2329, tmp_var);
      type_cast_2362_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2376_inst
    process(shr67_2373) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr67_2373, tmp_var);
      type_cast_2376_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2392_inst
    process(input_dim2x_x1_2319) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_2319, tmp_var);
      type_cast_2392_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2431_inst
    process(inc_2428) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2428, tmp_var);
      type_cast_2431_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2465_inst
    process(input_dim0x_x0_2462) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x0_2462, tmp_var);
      type_cast_2465_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_2138_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_2138_load_0_req_0;
      LOAD_padding_2138_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_2138_load_0_req_1;
      LOAD_padding_2138_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_2138_word_address_0;
      LOAD_padding_2138_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_2095_load_0 ptr_deref_2113_load_0 ptr_deref_2204_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_2095_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2113_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2204_load_0_req_0;
      ptr_deref_2095_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2113_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2204_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_2095_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2113_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2204_load_0_req_1;
      ptr_deref_2095_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2113_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2204_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2095_word_address_0 & ptr_deref_2113_word_address_0 & ptr_deref_2204_word_address_0;
      ptr_deref_2095_data_0 <= data_out(47 downto 32);
      ptr_deref_2113_data_0 <= data_out(31 downto 16);
      ptr_deref_2204_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 16,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(15 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_2123_load_0 ptr_deref_2148_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2123_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2148_load_0_req_0;
      ptr_deref_2123_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2148_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2123_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2148_load_0_req_1;
      ptr_deref_2123_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2148_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2123_word_address_0 & ptr_deref_2148_word_address_0;
      ptr_deref_2123_data_0 <= data_out(31 downto 16);
      ptr_deref_2148_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(15 downto 0),
          mtag => memory_space_8_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_2135_load_0 ptr_deref_2160_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2135_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2160_load_0_req_0;
      ptr_deref_2135_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2160_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2135_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2160_load_0_req_1;
      ptr_deref_2135_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2160_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2135_word_address_0 & ptr_deref_2160_word_address_0;
      ptr_deref_2135_data_0 <= data_out(31 downto 16);
      ptr_deref_2160_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(15 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_2172_load_0 ptr_deref_2184_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2172_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2184_load_0_req_0;
      ptr_deref_2172_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2184_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2172_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2184_load_0_req_1;
      ptr_deref_2172_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2184_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2172_word_address_0 & ptr_deref_2184_word_address_0;
      ptr_deref_2172_data_0 <= data_out(31 downto 16);
      ptr_deref_2184_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(15 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_2358_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2358_load_0_req_0;
      ptr_deref_2358_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2358_load_0_req_1;
      ptr_deref_2358_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2358_word_address_0;
      ptr_deref_2358_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(13 downto 0),
          mtag => memory_space_4_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(63 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_2387_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2387_store_0_req_0;
      ptr_deref_2387_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2387_store_0_req_1;
      ptr_deref_2387_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2387_word_address_0;
      data_in <= ptr_deref_2387_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(13 downto 0),
          mdata => memory_space_6_sr_data(63 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_2082_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_start_2082_inst_req_0;
      RPIPE_Block1_start_2082_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_start_2082_inst_req_1;
      RPIPE_Block1_start_2082_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_2083 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_2481_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_2481_inst_req_0;
      WPIPE_Block1_done_2481_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_2481_inst_req_1;
      WPIPE_Block1_done_2481_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_2083;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_7299_start: Boolean;
  signal convTransposeC_CP_7299_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block2_start_2491_inst_req_1 : boolean;
  signal ptr_deref_2522_load_0_req_1 : boolean;
  signal ptr_deref_2522_load_0_ack_1 : boolean;
  signal RPIPE_Block2_start_2491_inst_ack_1 : boolean;
  signal ptr_deref_2504_load_0_req_0 : boolean;
  signal ptr_deref_2504_load_0_ack_0 : boolean;
  signal ptr_deref_2544_load_0_ack_1 : boolean;
  signal ptr_deref_2544_load_0_req_1 : boolean;
  signal ptr_deref_2534_load_0_req_1 : boolean;
  signal ptr_deref_2534_load_0_ack_1 : boolean;
  signal ptr_deref_2544_load_0_req_0 : boolean;
  signal ptr_deref_2544_load_0_ack_0 : boolean;
  signal RPIPE_Block2_start_2491_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2491_inst_ack_0 : boolean;
  signal ptr_deref_2556_load_0_req_1 : boolean;
  signal ptr_deref_2556_load_0_req_0 : boolean;
  signal ptr_deref_2556_load_0_ack_0 : boolean;
  signal ptr_deref_2534_load_0_ack_0 : boolean;
  signal ptr_deref_2556_load_0_ack_1 : boolean;
  signal ptr_deref_2534_load_0_req_0 : boolean;
  signal ptr_deref_2522_load_0_ack_0 : boolean;
  signal ptr_deref_2522_load_0_req_0 : boolean;
  signal LOAD_padding_2559_load_0_ack_0 : boolean;
  signal ptr_deref_2504_load_0_ack_1 : boolean;
  signal ptr_deref_2504_load_0_req_1 : boolean;
  signal LOAD_padding_2559_load_0_req_1 : boolean;
  signal LOAD_padding_2559_load_0_ack_1 : boolean;
  signal LOAD_padding_2559_load_0_req_0 : boolean;
  signal ptr_deref_2569_load_0_req_0 : boolean;
  signal ptr_deref_2569_load_0_ack_0 : boolean;
  signal ptr_deref_2569_load_0_req_1 : boolean;
  signal ptr_deref_2569_load_0_ack_1 : boolean;
  signal ptr_deref_2581_load_0_req_0 : boolean;
  signal ptr_deref_2581_load_0_ack_0 : boolean;
  signal ptr_deref_2581_load_0_req_1 : boolean;
  signal ptr_deref_2581_load_0_ack_1 : boolean;
  signal ptr_deref_2593_load_0_req_0 : boolean;
  signal ptr_deref_2593_load_0_ack_0 : boolean;
  signal ptr_deref_2593_load_0_req_1 : boolean;
  signal ptr_deref_2593_load_0_ack_1 : boolean;
  signal ptr_deref_2605_load_0_req_0 : boolean;
  signal ptr_deref_2605_load_0_ack_0 : boolean;
  signal ptr_deref_2605_load_0_req_1 : boolean;
  signal ptr_deref_2605_load_0_ack_1 : boolean;
  signal type_cast_2609_inst_req_0 : boolean;
  signal type_cast_2609_inst_ack_0 : boolean;
  signal type_cast_2609_inst_req_1 : boolean;
  signal type_cast_2609_inst_ack_1 : boolean;
  signal type_cast_2613_inst_req_0 : boolean;
  signal type_cast_2613_inst_ack_0 : boolean;
  signal type_cast_2613_inst_req_1 : boolean;
  signal type_cast_2613_inst_ack_1 : boolean;
  signal type_cast_2623_inst_req_0 : boolean;
  signal type_cast_2623_inst_ack_0 : boolean;
  signal type_cast_2623_inst_req_1 : boolean;
  signal type_cast_2623_inst_ack_1 : boolean;
  signal type_cast_2742_inst_req_0 : boolean;
  signal type_cast_2742_inst_ack_0 : boolean;
  signal type_cast_2742_inst_req_1 : boolean;
  signal type_cast_2742_inst_ack_1 : boolean;
  signal type_cast_2756_inst_req_0 : boolean;
  signal type_cast_2756_inst_ack_0 : boolean;
  signal type_cast_2756_inst_req_1 : boolean;
  signal type_cast_2756_inst_ack_1 : boolean;
  signal array_obj_ref_2762_index_offset_req_0 : boolean;
  signal array_obj_ref_2762_index_offset_ack_0 : boolean;
  signal array_obj_ref_2762_index_offset_req_1 : boolean;
  signal array_obj_ref_2762_index_offset_ack_1 : boolean;
  signal addr_of_2763_final_reg_req_0 : boolean;
  signal addr_of_2763_final_reg_ack_0 : boolean;
  signal addr_of_2763_final_reg_req_1 : boolean;
  signal addr_of_2763_final_reg_ack_1 : boolean;
  signal ptr_deref_2767_load_0_req_0 : boolean;
  signal ptr_deref_2767_load_0_ack_0 : boolean;
  signal ptr_deref_2767_load_0_req_1 : boolean;
  signal ptr_deref_2767_load_0_ack_1 : boolean;
  signal type_cast_2772_inst_req_0 : boolean;
  signal type_cast_2772_inst_ack_0 : boolean;
  signal type_cast_2772_inst_req_1 : boolean;
  signal type_cast_2772_inst_ack_1 : boolean;
  signal type_cast_2786_inst_req_0 : boolean;
  signal type_cast_2786_inst_ack_0 : boolean;
  signal type_cast_2786_inst_req_1 : boolean;
  signal type_cast_2786_inst_ack_1 : boolean;
  signal array_obj_ref_2792_index_offset_req_0 : boolean;
  signal array_obj_ref_2792_index_offset_ack_0 : boolean;
  signal array_obj_ref_2792_index_offset_req_1 : boolean;
  signal array_obj_ref_2792_index_offset_ack_1 : boolean;
  signal addr_of_2793_final_reg_req_0 : boolean;
  signal addr_of_2793_final_reg_ack_0 : boolean;
  signal addr_of_2793_final_reg_req_1 : boolean;
  signal addr_of_2793_final_reg_ack_1 : boolean;
  signal ptr_deref_2796_store_0_req_0 : boolean;
  signal ptr_deref_2796_store_0_ack_0 : boolean;
  signal ptr_deref_2796_store_0_req_1 : boolean;
  signal ptr_deref_2796_store_0_ack_1 : boolean;
  signal type_cast_2802_inst_req_0 : boolean;
  signal type_cast_2802_inst_ack_0 : boolean;
  signal type_cast_2802_inst_req_1 : boolean;
  signal type_cast_2802_inst_ack_1 : boolean;
  signal if_stmt_2817_branch_req_0 : boolean;
  signal if_stmt_2817_branch_ack_1 : boolean;
  signal if_stmt_2817_branch_ack_0 : boolean;
  signal type_cast_2841_inst_req_0 : boolean;
  signal type_cast_2841_inst_ack_0 : boolean;
  signal type_cast_2841_inst_req_1 : boolean;
  signal type_cast_2841_inst_ack_1 : boolean;
  signal type_cast_2850_inst_req_0 : boolean;
  signal type_cast_2850_inst_ack_0 : boolean;
  signal type_cast_2850_inst_req_1 : boolean;
  signal type_cast_2850_inst_ack_1 : boolean;
  signal type_cast_2867_inst_req_0 : boolean;
  signal type_cast_2867_inst_ack_0 : boolean;
  signal type_cast_2867_inst_req_1 : boolean;
  signal type_cast_2867_inst_ack_1 : boolean;
  signal if_stmt_2874_branch_req_0 : boolean;
  signal if_stmt_2874_branch_ack_1 : boolean;
  signal if_stmt_2874_branch_ack_0 : boolean;
  signal WPIPE_Block2_done_2882_inst_req_0 : boolean;
  signal WPIPE_Block2_done_2882_inst_ack_0 : boolean;
  signal WPIPE_Block2_done_2882_inst_req_1 : boolean;
  signal WPIPE_Block2_done_2882_inst_ack_1 : boolean;
  signal phi_stmt_2649_req_0 : boolean;
  signal type_cast_2659_inst_req_0 : boolean;
  signal type_cast_2659_inst_ack_0 : boolean;
  signal type_cast_2659_inst_req_1 : boolean;
  signal type_cast_2659_inst_ack_1 : boolean;
  signal phi_stmt_2656_req_0 : boolean;
  signal type_cast_2655_inst_req_0 : boolean;
  signal type_cast_2655_inst_ack_0 : boolean;
  signal type_cast_2655_inst_req_1 : boolean;
  signal type_cast_2655_inst_ack_1 : boolean;
  signal phi_stmt_2649_req_1 : boolean;
  signal type_cast_2661_inst_req_0 : boolean;
  signal type_cast_2661_inst_ack_0 : boolean;
  signal type_cast_2661_inst_req_1 : boolean;
  signal type_cast_2661_inst_ack_1 : boolean;
  signal phi_stmt_2656_req_1 : boolean;
  signal phi_stmt_2649_ack_0 : boolean;
  signal phi_stmt_2656_ack_0 : boolean;
  signal type_cast_2721_inst_req_0 : boolean;
  signal type_cast_2721_inst_ack_0 : boolean;
  signal type_cast_2721_inst_req_1 : boolean;
  signal type_cast_2721_inst_ack_1 : boolean;
  signal phi_stmt_2715_req_1 : boolean;
  signal phi_stmt_2715_req_0 : boolean;
  signal phi_stmt_2715_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_7299_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_7299_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_7299_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_7299_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_7299: Block -- control-path 
    signal convTransposeC_CP_7299_elements: BooleanArray(87 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_7299_elements(0) <= convTransposeC_CP_7299_start;
    convTransposeC_CP_7299_symbol <= convTransposeC_CP_7299_elements(65);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_2489/branch_block_stmt_2489__entry__
      -- CP-element group 0: 	 branch_block_stmt_2489/assign_stmt_2492__entry__
      -- CP-element group 0: 	 branch_block_stmt_2489/$entry
      -- CP-element group 0: 	 branch_block_stmt_2489/assign_stmt_2492/$entry
      -- CP-element group 0: 	 branch_block_stmt_2489/assign_stmt_2492/RPIPE_Block2_start_2491_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2489/assign_stmt_2492/RPIPE_Block2_start_2491_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2489/assign_stmt_2492/RPIPE_Block2_start_2491_Sample/rr
      -- CP-element group 0: 	 $entry
      -- 
    rr_7347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(0), ack => RPIPE_Block2_start_2491_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2489/assign_stmt_2492/RPIPE_Block2_start_2491_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2489/assign_stmt_2492/RPIPE_Block2_start_2491_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_2489/assign_stmt_2492/RPIPE_Block2_start_2491_update_start_
      -- CP-element group 1: 	 branch_block_stmt_2489/assign_stmt_2492/RPIPE_Block2_start_2491_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_2489/assign_stmt_2492/RPIPE_Block2_start_2491_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_2489/assign_stmt_2492/RPIPE_Block2_start_2491_Update/$entry
      -- 
    ra_7348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2491_inst_ack_0, ack => convTransposeC_CP_7299_elements(1)); -- 
    cr_7352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(1), ack => RPIPE_Block2_start_2491_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	21 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	11 
    -- CP-element group 2:  members (262) 
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2492/RPIPE_Block2_start_2491_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646__entry__
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2492__exit__
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2492/RPIPE_Block2_start_2491_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2492/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2492/RPIPE_Block2_start_2491_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2609_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2609_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2609_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2613_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2613_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2613_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2623_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2623_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2623_Update/cr
      -- 
    ca_7353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2491_inst_ack_1, ack => convTransposeC_CP_7299_elements(2)); -- 
    cr_7450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => ptr_deref_2522_load_0_req_1); -- 
    rr_7389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => ptr_deref_2504_load_0_req_0); -- 
    cr_7550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => ptr_deref_2544_load_0_req_1); -- 
    cr_7500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => ptr_deref_2534_load_0_req_1); -- 
    rr_7539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => ptr_deref_2544_load_0_req_0); -- 
    cr_7600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => ptr_deref_2556_load_0_req_1); -- 
    rr_7589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => ptr_deref_2556_load_0_req_0); -- 
    rr_7489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => ptr_deref_2534_load_0_req_0); -- 
    rr_7439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => ptr_deref_2522_load_0_req_0); -- 
    cr_7400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => ptr_deref_2504_load_0_req_1); -- 
    cr_7633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => LOAD_padding_2559_load_0_req_1); -- 
    rr_7622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => LOAD_padding_2559_load_0_req_0); -- 
    rr_7672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => ptr_deref_2569_load_0_req_0); -- 
    cr_7683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => ptr_deref_2569_load_0_req_1); -- 
    rr_7722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => ptr_deref_2581_load_0_req_0); -- 
    cr_7733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => ptr_deref_2581_load_0_req_1); -- 
    rr_7772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => ptr_deref_2593_load_0_req_0); -- 
    cr_7783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => ptr_deref_2593_load_0_req_1); -- 
    rr_7822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => ptr_deref_2605_load_0_req_0); -- 
    cr_7833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => ptr_deref_2605_load_0_req_1); -- 
    cr_7852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => type_cast_2609_inst_req_1); -- 
    cr_7866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => type_cast_2613_inst_req_1); -- 
    cr_7880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(2), ack => type_cast_2623_inst_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_Sample/word_access_start/word_0/ra
      -- CP-element group 3: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_Sample/$exit
      -- 
    ra_7390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2504_load_0_ack_0, ack => convTransposeC_CP_7299_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	27 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_Update/ptr_deref_2504_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_Update/ptr_deref_2504_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_Update/ptr_deref_2504_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_Update/ptr_deref_2504_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2504_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2623_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2623_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2623_Sample/rr
      -- 
    ca_7401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2504_load_0_ack_1, ack => convTransposeC_CP_7299_elements(4)); -- 
    rr_7875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(4), ack => type_cast_2623_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_Sample/word_access_start/word_0/ra
      -- CP-element group 5: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_Sample/word_access_start/$exit
      -- 
    ra_7440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2522_load_0_ack_0, ack => convTransposeC_CP_7299_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	23 
    -- CP-element group 6:  members (12) 
      -- CP-element group 6: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_Update/ptr_deref_2522_Merge/merge_ack
      -- CP-element group 6: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_Update/ptr_deref_2522_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_Update/ptr_deref_2522_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_Update/ptr_deref_2522_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2609_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2522_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2609_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2609_Sample/rr
      -- 
    ca_7451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2522_load_0_ack_1, ack => convTransposeC_CP_7299_elements(6)); -- 
    rr_7847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(6), ack => type_cast_2609_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_Sample/word_access_start/word_0/ra
      -- 
    ra_7490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2534_load_0_ack_0, ack => convTransposeC_CP_7299_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	25 
    -- CP-element group 8:  members (12) 
      -- CP-element group 8: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_Update/ptr_deref_2534_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_Update/ptr_deref_2534_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_Update/ptr_deref_2534_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_Update/ptr_deref_2534_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2534_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2613_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2613_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2613_Sample/rr
      -- 
    ca_7501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2534_load_0_ack_1, ack => convTransposeC_CP_7299_elements(8)); -- 
    rr_7861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(8), ack => type_cast_2613_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_Sample/word_access_start/word_0/ra
      -- CP-element group 9: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_Sample/$exit
      -- 
    ra_7540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2544_load_0_ack_0, ack => convTransposeC_CP_7299_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	29 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_Update/ptr_deref_2544_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_Update/ptr_deref_2544_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_Update/ptr_deref_2544_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2544_Update/ptr_deref_2544_Merge/$entry
      -- 
    ca_7551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2544_load_0_ack_1, ack => convTransposeC_CP_7299_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_Sample/word_access_start/word_0/ra
      -- CP-element group 11: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_Sample/word_access_start/word_0/$exit
      -- 
    ra_7590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2556_load_0_ack_0, ack => convTransposeC_CP_7299_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	29 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_Update/ptr_deref_2556_Merge/merge_ack
      -- CP-element group 12: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_Update/ptr_deref_2556_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_Update/ptr_deref_2556_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_Update/ptr_deref_2556_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2556_update_completed_
      -- 
    ca_7601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2556_load_0_ack_1, ack => convTransposeC_CP_7299_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_Sample/word_access_start/word_0/ra
      -- CP-element group 13: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_Sample/word_access_start/word_0/$exit
      -- 
    ra_7623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2559_load_0_ack_0, ack => convTransposeC_CP_7299_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	29 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_Update/LOAD_padding_2559_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_Update/LOAD_padding_2559_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_Update/LOAD_padding_2559_Merge/merge_ack
      -- CP-element group 14: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/LOAD_padding_2559_Update/LOAD_padding_2559_Merge/$entry
      -- 
    ca_7634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2559_load_0_ack_1, ack => convTransposeC_CP_7299_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_Sample/word_access_start/word_0/ra
      -- 
    ra_7673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2569_load_0_ack_0, ack => convTransposeC_CP_7299_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	29 
    -- CP-element group 16:  members (9) 
      -- CP-element group 16: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_Update/ptr_deref_2569_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_Update/ptr_deref_2569_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_Update/ptr_deref_2569_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2569_Update/ptr_deref_2569_Merge/merge_ack
      -- 
    ca_7684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2569_load_0_ack_1, ack => convTransposeC_CP_7299_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_Sample/word_access_start/word_0/ra
      -- 
    ra_7723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2581_load_0_ack_0, ack => convTransposeC_CP_7299_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	29 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_Update/ptr_deref_2581_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_Update/ptr_deref_2581_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_Update/ptr_deref_2581_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2581_Update/ptr_deref_2581_Merge/merge_ack
      -- 
    ca_7734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2581_load_0_ack_1, ack => convTransposeC_CP_7299_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_Sample/word_access_start/word_0/ra
      -- 
    ra_7773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2593_load_0_ack_0, ack => convTransposeC_CP_7299_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	29 
    -- CP-element group 20:  members (9) 
      -- CP-element group 20: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_Update/ptr_deref_2593_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_Update/ptr_deref_2593_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_Update/ptr_deref_2593_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2593_Update/ptr_deref_2593_Merge/merge_ack
      -- 
    ca_7784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2593_load_0_ack_1, ack => convTransposeC_CP_7299_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	2 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_Sample/word_access_start/word_0/ra
      -- 
    ra_7823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2605_load_0_ack_0, ack => convTransposeC_CP_7299_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	29 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_Update/word_access_complete/word_0/ca
      -- CP-element group 22: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_Update/ptr_deref_2605_Merge/$entry
      -- CP-element group 22: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_Update/ptr_deref_2605_Merge/$exit
      -- CP-element group 22: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_Update/ptr_deref_2605_Merge/merge_req
      -- CP-element group 22: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/ptr_deref_2605_Update/ptr_deref_2605_Merge/merge_ack
      -- 
    ca_7834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2605_load_0_ack_1, ack => convTransposeC_CP_7299_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	6 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2609_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2609_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2609_Sample/ra
      -- 
    ra_7848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2609_inst_ack_0, ack => convTransposeC_CP_7299_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	29 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2609_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2609_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2609_Update/ca
      -- 
    ca_7853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2609_inst_ack_1, ack => convTransposeC_CP_7299_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	8 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2613_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2613_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2613_Sample/ra
      -- 
    ra_7862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2613_inst_ack_0, ack => convTransposeC_CP_7299_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2613_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2613_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2613_Update/ca
      -- 
    ca_7867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2613_inst_ack_1, ack => convTransposeC_CP_7299_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	4 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2623_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2623_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2623_Sample/ra
      -- 
    ra_7876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2623_inst_ack_0, ack => convTransposeC_CP_7299_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2623_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2623_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/type_cast_2623_Update/ca
      -- 
    ca_7881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2623_inst_ack_1, ack => convTransposeC_CP_7299_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  place  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: 	20 
    -- CP-element group 29: 	14 
    -- CP-element group 29: 	12 
    -- CP-element group 29: 	22 
    -- CP-element group 29: 	24 
    -- CP-element group 29: 	26 
    -- CP-element group 29: 	16 
    -- CP-element group 29: 	18 
    -- CP-element group 29: 	10 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	66 
    -- CP-element group 29: 	67 
    -- CP-element group 29: 	68 
    -- CP-element group 29:  members (14) 
      -- CP-element group 29: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter
      -- CP-element group 29: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646__exit__
      -- CP-element group 29: 	 branch_block_stmt_2489/assign_stmt_2501_to_assign_stmt_2646/$exit
      -- CP-element group 29: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 29: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/$entry
      -- CP-element group 29: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/$entry
      -- CP-element group 29: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2659/$entry
      -- CP-element group 29: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2659/SplitProtocol/$entry
      -- CP-element group 29: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2659/SplitProtocol/Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2659/SplitProtocol/Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2659/SplitProtocol/Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2659/SplitProtocol/Update/cr
      -- 
    rr_8279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(29), ack => type_cast_2659_inst_req_0); -- 
    cr_8284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(29), ack => type_cast_2659_inst_req_1); -- 
    convTransposeC_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeC_CP_7299_elements(28) & convTransposeC_CP_7299_elements(20) & convTransposeC_CP_7299_elements(14) & convTransposeC_CP_7299_elements(12) & convTransposeC_CP_7299_elements(22) & convTransposeC_CP_7299_elements(24) & convTransposeC_CP_7299_elements(26) & convTransposeC_CP_7299_elements(16) & convTransposeC_CP_7299_elements(18) & convTransposeC_CP_7299_elements(10);
      gj_convTransposeC_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_7299_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	87 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2742_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2742_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2742_Sample/ra
      -- 
    ra_7896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2742_inst_ack_0, ack => convTransposeC_CP_7299_elements(30)); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	87 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2742_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2742_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2742_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2756_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2756_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2756_Sample/rr
      -- 
    ca_7901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2742_inst_ack_1, ack => convTransposeC_CP_7299_elements(31)); -- 
    rr_7909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(31), ack => type_cast_2756_inst_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2756_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2756_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2756_Sample/ra
      -- 
    ra_7910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2756_inst_ack_0, ack => convTransposeC_CP_7299_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	87 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (16) 
      -- CP-element group 33: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2756_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2756_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2756_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_index_resized_1
      -- CP-element group 33: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_index_scaled_1
      -- CP-element group 33: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_index_computed_1
      -- CP-element group 33: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_index_resize_1/$entry
      -- CP-element group 33: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_index_resize_1/$exit
      -- CP-element group 33: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_index_resize_1/index_resize_req
      -- CP-element group 33: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_index_resize_1/index_resize_ack
      -- CP-element group 33: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_index_scale_1/$entry
      -- CP-element group 33: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_index_scale_1/$exit
      -- CP-element group 33: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_index_scale_1/scale_rename_req
      -- CP-element group 33: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_index_scale_1/scale_rename_ack
      -- CP-element group 33: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_final_index_sum_regn_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_final_index_sum_regn_Sample/req
      -- 
    ca_7915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2756_inst_ack_1, ack => convTransposeC_CP_7299_elements(33)); -- 
    req_7940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(33), ack => array_obj_ref_2762_index_offset_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	53 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_final_index_sum_regn_sample_complete
      -- CP-element group 34: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_final_index_sum_regn_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_final_index_sum_regn_Sample/ack
      -- 
    ack_7941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2762_index_offset_ack_0, ack => convTransposeC_CP_7299_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	87 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (11) 
      -- CP-element group 35: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2763_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_root_address_calculated
      -- CP-element group 35: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_offset_calculated
      -- CP-element group 35: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_final_index_sum_regn_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_final_index_sum_regn_Update/ack
      -- CP-element group 35: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_base_plus_offset/$entry
      -- CP-element group 35: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_base_plus_offset/$exit
      -- CP-element group 35: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_base_plus_offset/sum_rename_req
      -- CP-element group 35: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_base_plus_offset/sum_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2763_request/$entry
      -- CP-element group 35: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2763_request/req
      -- 
    ack_7946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2762_index_offset_ack_1, ack => convTransposeC_CP_7299_elements(35)); -- 
    req_7955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(35), ack => addr_of_2763_final_reg_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2763_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2763_request/$exit
      -- CP-element group 36: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2763_request/ack
      -- 
    ack_7956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2763_final_reg_ack_0, ack => convTransposeC_CP_7299_elements(36)); -- 
    -- CP-element group 37:  join  fork  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	87 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (24) 
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2763_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2763_complete/$exit
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2763_complete/ack
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_base_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_word_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_base_address_resized
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_base_addr_resize/$entry
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_base_addr_resize/$exit
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_base_addr_resize/base_resize_req
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_base_addr_resize/base_resize_ack
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_base_plus_offset/$entry
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_base_plus_offset/$exit
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_base_plus_offset/sum_rename_req
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_word_addrgen/$entry
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_word_addrgen/$exit
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_word_addrgen/root_register_req
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_word_addrgen/root_register_ack
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_Sample/word_access_start/$entry
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_Sample/word_access_start/word_0/$entry
      -- CP-element group 37: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_Sample/word_access_start/word_0/rr
      -- 
    ack_7961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2763_final_reg_ack_1, ack => convTransposeC_CP_7299_elements(37)); -- 
    rr_7994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(37), ack => ptr_deref_2767_load_0_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_Sample/word_access_start/$exit
      -- CP-element group 38: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_Sample/word_access_start/word_0/$exit
      -- CP-element group 38: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_Sample/word_access_start/word_0/ra
      -- 
    ra_7995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2767_load_0_ack_0, ack => convTransposeC_CP_7299_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	87 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	48 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_Update/word_access_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_Update/word_access_complete/word_0/$exit
      -- CP-element group 39: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_Update/word_access_complete/word_0/ca
      -- CP-element group 39: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_Update/ptr_deref_2767_Merge/$entry
      -- CP-element group 39: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_Update/ptr_deref_2767_Merge/$exit
      -- CP-element group 39: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_Update/ptr_deref_2767_Merge/merge_req
      -- CP-element group 39: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_Update/ptr_deref_2767_Merge/merge_ack
      -- 
    ca_8006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2767_load_0_ack_1, ack => convTransposeC_CP_7299_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	87 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2772_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2772_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2772_Sample/ra
      -- 
    ra_8020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2772_inst_ack_0, ack => convTransposeC_CP_7299_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	87 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2772_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2772_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2772_Update/ca
      -- CP-element group 41: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2786_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2786_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2786_Sample/rr
      -- 
    ca_8025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2772_inst_ack_1, ack => convTransposeC_CP_7299_elements(41)); -- 
    rr_8033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(41), ack => type_cast_2786_inst_req_0); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2786_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2786_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2786_Sample/ra
      -- 
    ra_8034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2786_inst_ack_0, ack => convTransposeC_CP_7299_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	87 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (16) 
      -- CP-element group 43: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2786_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2786_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2786_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_index_resized_1
      -- CP-element group 43: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_index_scaled_1
      -- CP-element group 43: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_index_computed_1
      -- CP-element group 43: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_index_resize_1/$entry
      -- CP-element group 43: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_index_resize_1/$exit
      -- CP-element group 43: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_index_resize_1/index_resize_req
      -- CP-element group 43: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_index_resize_1/index_resize_ack
      -- CP-element group 43: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_index_scale_1/$entry
      -- CP-element group 43: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_index_scale_1/$exit
      -- CP-element group 43: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_index_scale_1/scale_rename_req
      -- CP-element group 43: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_index_scale_1/scale_rename_ack
      -- CP-element group 43: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_final_index_sum_regn_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_final_index_sum_regn_Sample/req
      -- 
    ca_8039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2786_inst_ack_1, ack => convTransposeC_CP_7299_elements(43)); -- 
    req_8064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(43), ack => array_obj_ref_2792_index_offset_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	53 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_final_index_sum_regn_sample_complete
      -- CP-element group 44: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_final_index_sum_regn_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_final_index_sum_regn_Sample/ack
      -- 
    ack_8065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2792_index_offset_ack_0, ack => convTransposeC_CP_7299_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	87 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (11) 
      -- CP-element group 45: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2793_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_root_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_offset_calculated
      -- CP-element group 45: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_final_index_sum_regn_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_final_index_sum_regn_Update/ack
      -- CP-element group 45: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_base_plus_offset/$entry
      -- CP-element group 45: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_base_plus_offset/$exit
      -- CP-element group 45: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_base_plus_offset/sum_rename_req
      -- CP-element group 45: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_base_plus_offset/sum_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2793_request/$entry
      -- CP-element group 45: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2793_request/req
      -- 
    ack_8070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2792_index_offset_ack_1, ack => convTransposeC_CP_7299_elements(45)); -- 
    req_8079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(45), ack => addr_of_2793_final_reg_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2793_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2793_request/$exit
      -- CP-element group 46: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2793_request/ack
      -- 
    ack_8080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2793_final_reg_ack_0, ack => convTransposeC_CP_7299_elements(46)); -- 
    -- CP-element group 47:  fork  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	87 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (19) 
      -- CP-element group 47: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2793_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2793_complete/$exit
      -- CP-element group 47: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2793_complete/ack
      -- CP-element group 47: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_base_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_word_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_root_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_base_address_resized
      -- CP-element group 47: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_base_addr_resize/$entry
      -- CP-element group 47: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_base_addr_resize/$exit
      -- CP-element group 47: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_base_addr_resize/base_resize_req
      -- CP-element group 47: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_base_addr_resize/base_resize_ack
      -- CP-element group 47: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_base_plus_offset/$entry
      -- CP-element group 47: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_base_plus_offset/$exit
      -- CP-element group 47: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_base_plus_offset/sum_rename_req
      -- CP-element group 47: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_base_plus_offset/sum_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_word_addrgen/$entry
      -- CP-element group 47: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_word_addrgen/$exit
      -- CP-element group 47: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_word_addrgen/root_register_req
      -- CP-element group 47: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_word_addrgen/root_register_ack
      -- 
    ack_8085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2793_final_reg_ack_1, ack => convTransposeC_CP_7299_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: 	39 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (9) 
      -- CP-element group 48: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_Sample/ptr_deref_2796_Split/$entry
      -- CP-element group 48: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_Sample/ptr_deref_2796_Split/$exit
      -- CP-element group 48: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_Sample/ptr_deref_2796_Split/split_req
      -- CP-element group 48: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_Sample/ptr_deref_2796_Split/split_ack
      -- CP-element group 48: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_Sample/word_access_start/$entry
      -- CP-element group 48: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_Sample/word_access_start/word_0/$entry
      -- CP-element group 48: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_Sample/word_access_start/word_0/rr
      -- 
    rr_8123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(48), ack => ptr_deref_2796_store_0_req_0); -- 
    convTransposeC_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_7299_elements(47) & convTransposeC_CP_7299_elements(39);
      gj_convTransposeC_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_7299_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_Sample/word_access_start/$exit
      -- CP-element group 49: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_Sample/word_access_start/word_0/$exit
      -- CP-element group 49: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_Sample/word_access_start/word_0/ra
      -- 
    ra_8124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2796_store_0_ack_0, ack => convTransposeC_CP_7299_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	87 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_Update/word_access_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_Update/word_access_complete/word_0/$exit
      -- CP-element group 50: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_Update/word_access_complete/word_0/ca
      -- 
    ca_8135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2796_store_0_ack_1, ack => convTransposeC_CP_7299_elements(50)); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	87 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2802_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2802_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2802_Sample/ra
      -- 
    ra_8144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2802_inst_ack_0, ack => convTransposeC_CP_7299_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	87 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2802_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2802_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2802_Update/ca
      -- 
    ca_8149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2802_inst_ack_1, ack => convTransposeC_CP_7299_elements(52)); -- 
    -- CP-element group 53:  branch  join  transition  place  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: 	52 
    -- CP-element group 53: 	44 
    -- CP-element group 53: 	34 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (10) 
      -- CP-element group 53: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816__exit__
      -- CP-element group 53: 	 branch_block_stmt_2489/if_stmt_2817__entry__
      -- CP-element group 53: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/$exit
      -- CP-element group 53: 	 branch_block_stmt_2489/if_stmt_2817_dead_link/$entry
      -- CP-element group 53: 	 branch_block_stmt_2489/if_stmt_2817_eval_test/$entry
      -- CP-element group 53: 	 branch_block_stmt_2489/if_stmt_2817_eval_test/$exit
      -- CP-element group 53: 	 branch_block_stmt_2489/if_stmt_2817_eval_test/branch_req
      -- CP-element group 53: 	 branch_block_stmt_2489/R_cmp_2818_place
      -- CP-element group 53: 	 branch_block_stmt_2489/if_stmt_2817_if_link/$entry
      -- CP-element group 53: 	 branch_block_stmt_2489/if_stmt_2817_else_link/$entry
      -- 
    branch_req_8157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(53), ack => if_stmt_2817_branch_req_0); -- 
    convTransposeC_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_7299_elements(50) & convTransposeC_CP_7299_elements(52) & convTransposeC_CP_7299_elements(44) & convTransposeC_CP_7299_elements(34);
      gj_convTransposeC_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_7299_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	82 
    -- CP-element group 54: 	83 
    -- CP-element group 54:  members (24) 
      -- CP-element group 54: 	 branch_block_stmt_2489/assign_stmt_2829__entry__
      -- CP-element group 54: 	 branch_block_stmt_2489/assign_stmt_2829__exit__
      -- CP-element group 54: 	 branch_block_stmt_2489/ifx_xthen_whilex_xbody
      -- CP-element group 54: 	 branch_block_stmt_2489/merge_stmt_2823__exit__
      -- CP-element group 54: 	 branch_block_stmt_2489/if_stmt_2817_if_link/$exit
      -- CP-element group 54: 	 branch_block_stmt_2489/if_stmt_2817_if_link/if_choice_transition
      -- CP-element group 54: 	 branch_block_stmt_2489/whilex_xbody_ifx_xthen
      -- CP-element group 54: 	 branch_block_stmt_2489/assign_stmt_2829/$entry
      -- CP-element group 54: 	 branch_block_stmt_2489/assign_stmt_2829/$exit
      -- CP-element group 54: 	 branch_block_stmt_2489/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_2489/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2715/$entry
      -- CP-element group 54: 	 branch_block_stmt_2489/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/$entry
      -- CP-element group 54: 	 branch_block_stmt_2489/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/$entry
      -- CP-element group 54: 	 branch_block_stmt_2489/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/SplitProtocol/$entry
      -- CP-element group 54: 	 branch_block_stmt_2489/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/SplitProtocol/Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_2489/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/SplitProtocol/Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_2489/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/SplitProtocol/Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_2489/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/SplitProtocol/Update/cr
      -- CP-element group 54: 	 branch_block_stmt_2489/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_2489/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 54: 	 branch_block_stmt_2489/merge_stmt_2823_PhiReqMerge
      -- CP-element group 54: 	 branch_block_stmt_2489/merge_stmt_2823_PhiAck/$entry
      -- CP-element group 54: 	 branch_block_stmt_2489/merge_stmt_2823_PhiAck/$exit
      -- CP-element group 54: 	 branch_block_stmt_2489/merge_stmt_2823_PhiAck/dummy
      -- 
    if_choice_transition_8162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2817_branch_ack_1, ack => convTransposeC_CP_7299_elements(54)); -- 
    rr_8360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(54), ack => type_cast_2721_inst_req_0); -- 
    cr_8365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(54), ack => type_cast_2721_inst_req_1); -- 
    -- CP-element group 55:  fork  transition  place  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	59 
    -- CP-element group 55: 	61 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_2489/merge_stmt_2831__exit__
      -- CP-element group 55: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873__entry__
      -- CP-element group 55: 	 branch_block_stmt_2489/if_stmt_2817_else_link/$exit
      -- CP-element group 55: 	 branch_block_stmt_2489/if_stmt_2817_else_link/else_choice_transition
      -- CP-element group 55: 	 branch_block_stmt_2489/whilex_xbody_ifx_xelse
      -- CP-element group 55: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/$entry
      -- CP-element group 55: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2841_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2841_update_start_
      -- CP-element group 55: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2841_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2841_Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2841_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2841_Update/cr
      -- CP-element group 55: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2850_update_start_
      -- CP-element group 55: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2850_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2850_Update/cr
      -- CP-element group 55: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2867_update_start_
      -- CP-element group 55: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2867_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2867_Update/cr
      -- CP-element group 55: 	 branch_block_stmt_2489/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 55: 	 branch_block_stmt_2489/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 55: 	 branch_block_stmt_2489/merge_stmt_2831_PhiReqMerge
      -- CP-element group 55: 	 branch_block_stmt_2489/merge_stmt_2831_PhiAck/$entry
      -- CP-element group 55: 	 branch_block_stmt_2489/merge_stmt_2831_PhiAck/$exit
      -- CP-element group 55: 	 branch_block_stmt_2489/merge_stmt_2831_PhiAck/dummy
      -- 
    else_choice_transition_8166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2817_branch_ack_0, ack => convTransposeC_CP_7299_elements(55)); -- 
    rr_8182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(55), ack => type_cast_2841_inst_req_0); -- 
    cr_8187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(55), ack => type_cast_2841_inst_req_1); -- 
    cr_8201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(55), ack => type_cast_2850_inst_req_1); -- 
    cr_8215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(55), ack => type_cast_2867_inst_req_1); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2841_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2841_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2841_Sample/ra
      -- 
    ra_8183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2841_inst_ack_0, ack => convTransposeC_CP_7299_elements(56)); -- 
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2841_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2841_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2841_Update/ca
      -- CP-element group 57: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2850_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2850_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2850_Sample/rr
      -- 
    ca_8188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2841_inst_ack_1, ack => convTransposeC_CP_7299_elements(57)); -- 
    rr_8196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(57), ack => type_cast_2850_inst_req_0); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2850_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2850_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2850_Sample/ra
      -- 
    ra_8197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2850_inst_ack_0, ack => convTransposeC_CP_7299_elements(58)); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	55 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2850_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2850_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2850_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2867_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2867_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2867_Sample/rr
      -- 
    ca_8202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2850_inst_ack_1, ack => convTransposeC_CP_7299_elements(59)); -- 
    rr_8210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(59), ack => type_cast_2867_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2867_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2867_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2867_Sample/ra
      -- 
    ra_8211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2867_inst_ack_0, ack => convTransposeC_CP_7299_elements(60)); -- 
    -- CP-element group 61:  branch  transition  place  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	55 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (13) 
      -- CP-element group 61: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873__exit__
      -- CP-element group 61: 	 branch_block_stmt_2489/if_stmt_2874__entry__
      -- CP-element group 61: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/$exit
      -- CP-element group 61: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2867_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2867_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_2489/assign_stmt_2837_to_assign_stmt_2873/type_cast_2867_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_2489/if_stmt_2874_dead_link/$entry
      -- CP-element group 61: 	 branch_block_stmt_2489/if_stmt_2874_eval_test/$entry
      -- CP-element group 61: 	 branch_block_stmt_2489/if_stmt_2874_eval_test/$exit
      -- CP-element group 61: 	 branch_block_stmt_2489/if_stmt_2874_eval_test/branch_req
      -- CP-element group 61: 	 branch_block_stmt_2489/R_cmp97_2875_place
      -- CP-element group 61: 	 branch_block_stmt_2489/if_stmt_2874_if_link/$entry
      -- CP-element group 61: 	 branch_block_stmt_2489/if_stmt_2874_else_link/$entry
      -- 
    ca_8216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2867_inst_ack_1, ack => convTransposeC_CP_7299_elements(61)); -- 
    branch_req_8224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(61), ack => if_stmt_2874_branch_req_0); -- 
    -- CP-element group 62:  merge  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (15) 
      -- CP-element group 62: 	 branch_block_stmt_2489/merge_stmt_2880__exit__
      -- CP-element group 62: 	 branch_block_stmt_2489/assign_stmt_2884__entry__
      -- CP-element group 62: 	 branch_block_stmt_2489/if_stmt_2874_if_link/$exit
      -- CP-element group 62: 	 branch_block_stmt_2489/if_stmt_2874_if_link/if_choice_transition
      -- CP-element group 62: 	 branch_block_stmt_2489/ifx_xelse_whilex_xend
      -- CP-element group 62: 	 branch_block_stmt_2489/assign_stmt_2884/$entry
      -- CP-element group 62: 	 branch_block_stmt_2489/assign_stmt_2884/WPIPE_Block2_done_2882_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_2489/assign_stmt_2884/WPIPE_Block2_done_2882_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_2489/assign_stmt_2884/WPIPE_Block2_done_2882_Sample/req
      -- CP-element group 62: 	 branch_block_stmt_2489/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 62: 	 branch_block_stmt_2489/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 62: 	 branch_block_stmt_2489/merge_stmt_2880_PhiReqMerge
      -- CP-element group 62: 	 branch_block_stmt_2489/merge_stmt_2880_PhiAck/$entry
      -- CP-element group 62: 	 branch_block_stmt_2489/merge_stmt_2880_PhiAck/$exit
      -- CP-element group 62: 	 branch_block_stmt_2489/merge_stmt_2880_PhiAck/dummy
      -- 
    if_choice_transition_8229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2874_branch_ack_1, ack => convTransposeC_CP_7299_elements(62)); -- 
    req_8246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(62), ack => WPIPE_Block2_done_2882_inst_req_0); -- 
    -- CP-element group 63:  fork  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	72 
    -- CP-element group 63: 	71 
    -- CP-element group 63: 	74 
    -- CP-element group 63: 	75 
    -- CP-element group 63:  members (20) 
      -- CP-element group 63: 	 branch_block_stmt_2489/if_stmt_2874_else_link/$exit
      -- CP-element group 63: 	 branch_block_stmt_2489/if_stmt_2874_else_link/else_choice_transition
      -- CP-element group 63: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 63: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 63: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/$entry
      -- CP-element group 63: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/$entry
      -- CP-element group 63: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/$entry
      -- CP-element group 63: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/SplitProtocol/$entry
      -- CP-element group 63: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/SplitProtocol/Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/SplitProtocol/Sample/rr
      -- CP-element group 63: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/SplitProtocol/Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/SplitProtocol/Update/cr
      -- CP-element group 63: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/$entry
      -- CP-element group 63: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/$entry
      -- CP-element group 63: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2661/$entry
      -- CP-element group 63: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2661/SplitProtocol/$entry
      -- CP-element group 63: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2661/SplitProtocol/Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2661/SplitProtocol/Sample/rr
      -- CP-element group 63: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2661/SplitProtocol/Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2661/SplitProtocol/Update/cr
      -- 
    else_choice_transition_8233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2874_branch_ack_0, ack => convTransposeC_CP_7299_elements(63)); -- 
    rr_8305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(63), ack => type_cast_2655_inst_req_0); -- 
    cr_8310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(63), ack => type_cast_2655_inst_req_1); -- 
    rr_8328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(63), ack => type_cast_2661_inst_req_0); -- 
    cr_8333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(63), ack => type_cast_2661_inst_req_1); -- 
    -- CP-element group 64:  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (6) 
      -- CP-element group 64: 	 branch_block_stmt_2489/assign_stmt_2884/WPIPE_Block2_done_2882_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2489/assign_stmt_2884/WPIPE_Block2_done_2882_update_start_
      -- CP-element group 64: 	 branch_block_stmt_2489/assign_stmt_2884/WPIPE_Block2_done_2882_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2489/assign_stmt_2884/WPIPE_Block2_done_2882_Sample/ack
      -- CP-element group 64: 	 branch_block_stmt_2489/assign_stmt_2884/WPIPE_Block2_done_2882_Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_2489/assign_stmt_2884/WPIPE_Block2_done_2882_Update/req
      -- 
    ack_8247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2882_inst_ack_0, ack => convTransposeC_CP_7299_elements(64)); -- 
    req_8251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(64), ack => WPIPE_Block2_done_2882_inst_req_1); -- 
    -- CP-element group 65:  transition  place  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (16) 
      -- CP-element group 65: 	 $exit
      -- CP-element group 65: 	 branch_block_stmt_2489/branch_block_stmt_2489__exit__
      -- CP-element group 65: 	 branch_block_stmt_2489/assign_stmt_2884__exit__
      -- CP-element group 65: 	 branch_block_stmt_2489/$exit
      -- CP-element group 65: 	 branch_block_stmt_2489/return__
      -- CP-element group 65: 	 branch_block_stmt_2489/merge_stmt_2886__exit__
      -- CP-element group 65: 	 branch_block_stmt_2489/assign_stmt_2884/$exit
      -- CP-element group 65: 	 branch_block_stmt_2489/assign_stmt_2884/WPIPE_Block2_done_2882_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2489/assign_stmt_2884/WPIPE_Block2_done_2882_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2489/assign_stmt_2884/WPIPE_Block2_done_2882_Update/ack
      -- CP-element group 65: 	 branch_block_stmt_2489/return___PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_2489/return___PhiReq/$exit
      -- CP-element group 65: 	 branch_block_stmt_2489/merge_stmt_2886_PhiReqMerge
      -- CP-element group 65: 	 branch_block_stmt_2489/merge_stmt_2886_PhiAck/$entry
      -- CP-element group 65: 	 branch_block_stmt_2489/merge_stmt_2886_PhiAck/$exit
      -- CP-element group 65: 	 branch_block_stmt_2489/merge_stmt_2886_PhiAck/dummy
      -- 
    ack_8252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2882_inst_ack_1, ack => convTransposeC_CP_7299_elements(65)); -- 
    -- CP-element group 66:  transition  output  delay-element  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	29 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	70 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/$exit
      -- CP-element group 66: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/$exit
      -- CP-element group 66: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2653_konst_delay_trans
      -- CP-element group 66: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/phi_stmt_2649_req
      -- 
    phi_stmt_2649_req_8263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2649_req_8263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(66), ack => phi_stmt_2649_req_0); -- 
    -- Element group convTransposeC_CP_7299_elements(66) is a control-delay.
    cp_element_66_delay: control_delay_element  generic map(name => " 66_delay", delay_value => 1)  port map(req => convTransposeC_CP_7299_elements(29), ack => convTransposeC_CP_7299_elements(66), clk => clk, reset =>reset);
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	29 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2659/SplitProtocol/Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2659/SplitProtocol/Sample/ra
      -- 
    ra_8280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2659_inst_ack_0, ack => convTransposeC_CP_7299_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	29 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2659/SplitProtocol/Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2659/SplitProtocol/Update/ca
      -- 
    ca_8285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2659_inst_ack_1, ack => convTransposeC_CP_7299_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (5) 
      -- CP-element group 69: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/$exit
      -- CP-element group 69: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/$exit
      -- CP-element group 69: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2659/$exit
      -- CP-element group 69: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2659/SplitProtocol/$exit
      -- CP-element group 69: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_req
      -- 
    phi_stmt_2656_req_8286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2656_req_8286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(69), ack => phi_stmt_2656_req_0); -- 
    convTransposeC_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_7299_elements(67) & convTransposeC_CP_7299_elements(68);
      gj_convTransposeC_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_7299_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  join  transition  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	66 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	78 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_2489/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_7299_elements(66) & convTransposeC_CP_7299_elements(69);
      gj_convTransposeC_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_7299_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	63 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/SplitProtocol/Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/SplitProtocol/Sample/ra
      -- 
    ra_8306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2655_inst_ack_0, ack => convTransposeC_CP_7299_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	63 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/SplitProtocol/Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/SplitProtocol/Update/ca
      -- 
    ca_8311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2655_inst_ack_1, ack => convTransposeC_CP_7299_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	77 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/$exit
      -- CP-element group 73: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/$exit
      -- CP-element group 73: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/$exit
      -- CP-element group 73: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/SplitProtocol/$exit
      -- CP-element group 73: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2649/phi_stmt_2649_req
      -- 
    phi_stmt_2649_req_8312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2649_req_8312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(73), ack => phi_stmt_2649_req_1); -- 
    convTransposeC_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_7299_elements(72) & convTransposeC_CP_7299_elements(71);
      gj_convTransposeC_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_7299_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	63 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2661/SplitProtocol/Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2661/SplitProtocol/Sample/ra
      -- 
    ra_8329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2661_inst_ack_0, ack => convTransposeC_CP_7299_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	63 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2661/SplitProtocol/Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2661/SplitProtocol/Update/ca
      -- 
    ca_8334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2661_inst_ack_1, ack => convTransposeC_CP_7299_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/$exit
      -- CP-element group 76: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2661/$exit
      -- CP-element group 76: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_sources/type_cast_2661/SplitProtocol/$exit
      -- CP-element group 76: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2656/phi_stmt_2656_req
      -- 
    phi_stmt_2656_req_8335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2656_req_8335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(76), ack => phi_stmt_2656_req_1); -- 
    convTransposeC_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_7299_elements(74) & convTransposeC_CP_7299_elements(75);
      gj_convTransposeC_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_7299_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	73 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_2489/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_7299_elements(73) & convTransposeC_CP_7299_elements(76);
      gj_convTransposeC_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_7299_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  merge  fork  transition  place  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	70 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2489/merge_stmt_2648_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_2489/merge_stmt_2648_PhiAck/$entry
      -- 
    convTransposeC_CP_7299_elements(78) <= OrReduce(convTransposeC_CP_7299_elements(70) & convTransposeC_CP_7299_elements(77));
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_2489/merge_stmt_2648_PhiAck/phi_stmt_2649_ack
      -- 
    phi_stmt_2649_ack_8340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2649_ack_0, ack => convTransposeC_CP_7299_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_2489/merge_stmt_2648_PhiAck/phi_stmt_2656_ack
      -- 
    phi_stmt_2656_ack_8341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2656_ack_0, ack => convTransposeC_CP_7299_elements(80)); -- 
    -- CP-element group 81:  join  transition  place  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (10) 
      -- CP-element group 81: 	 branch_block_stmt_2489/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 81: 	 branch_block_stmt_2489/merge_stmt_2648__exit__
      -- CP-element group 81: 	 branch_block_stmt_2489/assign_stmt_2667_to_assign_stmt_2712__entry__
      -- CP-element group 81: 	 branch_block_stmt_2489/assign_stmt_2667_to_assign_stmt_2712__exit__
      -- CP-element group 81: 	 branch_block_stmt_2489/assign_stmt_2667_to_assign_stmt_2712/$entry
      -- CP-element group 81: 	 branch_block_stmt_2489/assign_stmt_2667_to_assign_stmt_2712/$exit
      -- CP-element group 81: 	 branch_block_stmt_2489/merge_stmt_2648_PhiAck/$exit
      -- CP-element group 81: 	 branch_block_stmt_2489/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 81: 	 branch_block_stmt_2489/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2715/$entry
      -- CP-element group 81: 	 branch_block_stmt_2489/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/$entry
      -- 
    convTransposeC_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_7299_elements(79) & convTransposeC_CP_7299_elements(80);
      gj_convTransposeC_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_7299_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	54 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2489/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2489/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/SplitProtocol/Sample/ra
      -- 
    ra_8361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2721_inst_ack_0, ack => convTransposeC_CP_7299_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	54 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2489/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2489/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/SplitProtocol/Update/ca
      -- 
    ca_8366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2721_inst_ack_1, ack => convTransposeC_CP_7299_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (6) 
      -- CP-element group 84: 	 branch_block_stmt_2489/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 84: 	 branch_block_stmt_2489/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2715/$exit
      -- CP-element group 84: 	 branch_block_stmt_2489/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2489/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/$exit
      -- CP-element group 84: 	 branch_block_stmt_2489/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2721/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2489/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_req
      -- 
    phi_stmt_2715_req_8367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2715_req_8367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(84), ack => phi_stmt_2715_req_1); -- 
    convTransposeC_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_7299_elements(82) & convTransposeC_CP_7299_elements(83);
      gj_convTransposeC_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_7299_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  output  delay-element  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	81 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (5) 
      -- CP-element group 85: 	 branch_block_stmt_2489/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 85: 	 branch_block_stmt_2489/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2715/$exit
      -- CP-element group 85: 	 branch_block_stmt_2489/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/$exit
      -- CP-element group 85: 	 branch_block_stmt_2489/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_sources/type_cast_2719_konst_delay_trans
      -- CP-element group 85: 	 branch_block_stmt_2489/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2715/phi_stmt_2715_req
      -- 
    phi_stmt_2715_req_8378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2715_req_8378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(85), ack => phi_stmt_2715_req_0); -- 
    -- Element group convTransposeC_CP_7299_elements(85) is a control-delay.
    cp_element_85_delay: control_delay_element  generic map(name => " 85_delay", delay_value => 1)  port map(req => convTransposeC_CP_7299_elements(81), ack => convTransposeC_CP_7299_elements(85), clk => clk, reset =>reset);
    -- CP-element group 86:  merge  transition  place  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2489/merge_stmt_2714_PhiReqMerge
      -- CP-element group 86: 	 branch_block_stmt_2489/merge_stmt_2714_PhiAck/$entry
      -- 
    convTransposeC_CP_7299_elements(86) <= OrReduce(convTransposeC_CP_7299_elements(85) & convTransposeC_CP_7299_elements(84));
    -- CP-element group 87:  fork  transition  place  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	41 
    -- CP-element group 87: 	43 
    -- CP-element group 87: 	47 
    -- CP-element group 87: 	45 
    -- CP-element group 87: 	50 
    -- CP-element group 87: 	51 
    -- CP-element group 87: 	40 
    -- CP-element group 87: 	52 
    -- CP-element group 87: 	30 
    -- CP-element group 87: 	31 
    -- CP-element group 87: 	33 
    -- CP-element group 87: 	35 
    -- CP-element group 87: 	37 
    -- CP-element group 87: 	39 
    -- CP-element group 87:  members (51) 
      -- CP-element group 87: 	 branch_block_stmt_2489/merge_stmt_2714__exit__
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816__entry__
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/$entry
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2742_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2742_update_start_
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2742_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2742_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2742_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2742_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2756_update_start_
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2756_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2756_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2763_update_start_
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_final_index_sum_regn_update_start
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_final_index_sum_regn_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2762_final_index_sum_regn_Update/req
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2763_complete/$entry
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2763_complete/req
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_update_start_
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_Update/word_access_complete/$entry
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_Update/word_access_complete/word_0/$entry
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2767_Update/word_access_complete/word_0/cr
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2772_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2772_update_start_
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2772_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2772_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2772_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2772_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2786_update_start_
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2786_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2786_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2793_update_start_
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_final_index_sum_regn_update_start
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_final_index_sum_regn_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/array_obj_ref_2792_final_index_sum_regn_Update/req
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2793_complete/$entry
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/addr_of_2793_complete/req
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_update_start_
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_Update/word_access_complete/$entry
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_Update/word_access_complete/word_0/$entry
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/ptr_deref_2796_Update/word_access_complete/word_0/cr
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2802_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2802_update_start_
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2802_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2802_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2802_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_2489/assign_stmt_2728_to_assign_stmt_2816/type_cast_2802_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_2489/merge_stmt_2714_PhiAck/$exit
      -- CP-element group 87: 	 branch_block_stmt_2489/merge_stmt_2714_PhiAck/phi_stmt_2715_ack
      -- 
    phi_stmt_2715_ack_8383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2715_ack_0, ack => convTransposeC_CP_7299_elements(87)); -- 
    rr_7895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(87), ack => type_cast_2742_inst_req_0); -- 
    cr_7900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(87), ack => type_cast_2742_inst_req_1); -- 
    cr_7914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(87), ack => type_cast_2756_inst_req_1); -- 
    req_7945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(87), ack => array_obj_ref_2762_index_offset_req_1); -- 
    req_7960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(87), ack => addr_of_2763_final_reg_req_1); -- 
    cr_8005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(87), ack => ptr_deref_2767_load_0_req_1); -- 
    rr_8019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(87), ack => type_cast_2772_inst_req_0); -- 
    cr_8024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(87), ack => type_cast_2772_inst_req_1); -- 
    cr_8038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(87), ack => type_cast_2786_inst_req_1); -- 
    req_8069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(87), ack => array_obj_ref_2792_index_offset_req_1); -- 
    req_8084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(87), ack => addr_of_2793_final_reg_req_1); -- 
    cr_8134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(87), ack => ptr_deref_2796_store_0_req_1); -- 
    rr_8143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(87), ack => type_cast_2802_inst_req_0); -- 
    cr_8148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_7299_elements(87), ack => type_cast_2802_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2750_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2780_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_2559_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_2559_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom69_2791_resized : std_logic_vector(13 downto 0);
    signal R_idxprom69_2791_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2761_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2761_scaled : std_logic_vector(13 downto 0);
    signal add21_2733 : std_logic_vector(15 downto 0);
    signal add61_2738 : std_logic_vector(15 downto 0);
    signal add74_2809 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2762_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2762_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2762_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2762_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2762_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2762_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2792_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2792_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2792_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2792_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2792_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2792_root_address : std_logic_vector(13 downto 0);
    signal arrayidx70_2794 : std_logic_vector(31 downto 0);
    signal arrayidx_2764 : std_logic_vector(31 downto 0);
    signal call_2492 : std_logic_vector(15 downto 0);
    signal cmp88_2847 : std_logic_vector(0 downto 0);
    signal cmp97_2873 : std_logic_vector(0 downto 0);
    signal cmp_2816 : std_logic_vector(0 downto 0);
    signal conv64_2743 : std_logic_vector(31 downto 0);
    signal conv67_2773 : std_logic_vector(31 downto 0);
    signal conv73_2803 : std_logic_vector(31 downto 0);
    signal conv76_2610 : std_logic_vector(31 downto 0);
    signal conv84_2842 : std_logic_vector(31 downto 0);
    signal conv86_2614 : std_logic_vector(31 downto 0);
    signal conv94_2868 : std_logic_vector(31 downto 0);
    signal conv96_2624 : std_logic_vector(31 downto 0);
    signal div87_2620 : std_logic_vector(31 downto 0);
    signal div_2511 : std_logic_vector(15 downto 0);
    signal iNsTr_10_2602 : std_logic_vector(31 downto 0);
    signal iNsTr_2_2501 : std_logic_vector(31 downto 0);
    signal iNsTr_3_2519 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2531 : std_logic_vector(31 downto 0);
    signal iNsTr_5_2541 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2553 : std_logic_vector(31 downto 0);
    signal iNsTr_7_2566 : std_logic_vector(31 downto 0);
    signal iNsTr_8_2578 : std_logic_vector(31 downto 0);
    signal iNsTr_9_2590 : std_logic_vector(31 downto 0);
    signal idxprom69_2787 : std_logic_vector(63 downto 0);
    signal idxprom_2757 : std_logic_vector(63 downto 0);
    signal inc92_2851 : std_logic_vector(15 downto 0);
    signal inc92x_xinput_dim0x_x2_2856 : std_logic_vector(15 downto 0);
    signal inc_2837 : std_logic_vector(15 downto 0);
    signal indvar_2715 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2829 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2656 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2649 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2863 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2728 : std_logic_vector(15 downto 0);
    signal ptr_deref_2504_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2504_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2504_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2504_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2504_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2522_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2522_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2522_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2522_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2522_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2534_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2534_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2534_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2534_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2534_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2544_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2544_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2544_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2544_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2544_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2556_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2556_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2556_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2556_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2556_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2569_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2569_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2569_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2569_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2569_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2581_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2581_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2581_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2581_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2581_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2593_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2593_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2593_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2593_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2593_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2605_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2605_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2605_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2605_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2605_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2767_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2767_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2767_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2767_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2767_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2796_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2796_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2796_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2796_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2796_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2796_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr68_2782 : std_logic_vector(31 downto 0);
    signal shr_2752 : std_logic_vector(31 downto 0);
    signal tmp10_2697 : std_logic_vector(15 downto 0);
    signal tmp11_2702 : std_logic_vector(15 downto 0);
    signal tmp125_2667 : std_logic_vector(15 downto 0);
    signal tmp126_2672 : std_logic_vector(15 downto 0);
    signal tmp127_2677 : std_logic_vector(15 downto 0);
    signal tmp12_2523 : std_logic_vector(15 downto 0);
    signal tmp13_2707 : std_logic_vector(15 downto 0);
    signal tmp14_2712 : std_logic_vector(15 downto 0);
    signal tmp16_2535 : std_logic_vector(15 downto 0);
    signal tmp25_2545 : std_logic_vector(15 downto 0);
    signal tmp28_2557 : std_logic_vector(15 downto 0);
    signal tmp31_2560 : std_logic_vector(15 downto 0);
    signal tmp37_2570 : std_logic_vector(15 downto 0);
    signal tmp3_2630 : std_logic_vector(15 downto 0);
    signal tmp40_2582 : std_logic_vector(15 downto 0);
    signal tmp4_2635 : std_logic_vector(15 downto 0);
    signal tmp50_2594 : std_logic_vector(15 downto 0);
    signal tmp54_2606 : std_logic_vector(15 downto 0);
    signal tmp5_2682 : std_logic_vector(15 downto 0);
    signal tmp65_2768 : std_logic_vector(63 downto 0);
    signal tmp6_2687 : std_logic_vector(15 downto 0);
    signal tmp7_2641 : std_logic_vector(15 downto 0);
    signal tmp8_2646 : std_logic_vector(15 downto 0);
    signal tmp9_2692 : std_logic_vector(15 downto 0);
    signal tmp_2505 : std_logic_vector(15 downto 0);
    signal type_cast_2509_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2618_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2628_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2639_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2653_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2655_wire : std_logic_vector(15 downto 0);
    signal type_cast_2659_wire : std_logic_vector(15 downto 0);
    signal type_cast_2661_wire : std_logic_vector(15 downto 0);
    signal type_cast_2719_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2721_wire : std_logic_vector(15 downto 0);
    signal type_cast_2726_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2741_wire : std_logic_vector(31 downto 0);
    signal type_cast_2746_wire : std_logic_vector(31 downto 0);
    signal type_cast_2749_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2755_wire : std_logic_vector(63 downto 0);
    signal type_cast_2771_wire : std_logic_vector(31 downto 0);
    signal type_cast_2776_wire : std_logic_vector(31 downto 0);
    signal type_cast_2779_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2785_wire : std_logic_vector(63 downto 0);
    signal type_cast_2801_wire : std_logic_vector(31 downto 0);
    signal type_cast_2807_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2812_wire : std_logic_vector(31 downto 0);
    signal type_cast_2814_wire : std_logic_vector(31 downto 0);
    signal type_cast_2827_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2835_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2840_wire : std_logic_vector(31 downto 0);
    signal type_cast_2860_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2866_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_2559_word_address_0 <= "0";
    array_obj_ref_2762_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2762_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2762_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2762_resized_base_address <= "00000000000000";
    array_obj_ref_2792_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2792_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2792_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2792_resized_base_address <= "00000000000000";
    iNsTr_10_2602 <= "00000000000000000000000000000101";
    iNsTr_2_2501 <= "00000000000000000000000000000100";
    iNsTr_3_2519 <= "00000000000000000000000000000110";
    iNsTr_4_2531 <= "00000000000000000000000000000101";
    iNsTr_5_2541 <= "00000000000000000000000000000000";
    iNsTr_6_2553 <= "00000000000000000000000000000101";
    iNsTr_7_2566 <= "00000000000000000000000000000001";
    iNsTr_8_2578 <= "00000000000000000000000000000110";
    iNsTr_9_2590 <= "00000000000000000000000000000110";
    ptr_deref_2504_word_offset_0 <= "0000000";
    ptr_deref_2522_word_offset_0 <= "0000000";
    ptr_deref_2534_word_offset_0 <= "0000000";
    ptr_deref_2544_word_offset_0 <= "0";
    ptr_deref_2556_word_offset_0 <= "0000000";
    ptr_deref_2569_word_offset_0 <= "0";
    ptr_deref_2581_word_offset_0 <= "0000000";
    ptr_deref_2593_word_offset_0 <= "0000000";
    ptr_deref_2605_word_offset_0 <= "0000000";
    ptr_deref_2767_word_offset_0 <= "00000000000000";
    ptr_deref_2796_word_offset_0 <= "00000000000000";
    type_cast_2509_wire_constant <= "0000000000000001";
    type_cast_2618_wire_constant <= "00000000000000000000000000000001";
    type_cast_2628_wire_constant <= "1111111111111111";
    type_cast_2639_wire_constant <= "1111111111111111";
    type_cast_2653_wire_constant <= "0000000000000000";
    type_cast_2719_wire_constant <= "0000000000000000";
    type_cast_2726_wire_constant <= "0000000000000100";
    type_cast_2749_wire_constant <= "00000000000000000000000000000010";
    type_cast_2779_wire_constant <= "00000000000000000000000000000010";
    type_cast_2807_wire_constant <= "00000000000000000000000000000100";
    type_cast_2827_wire_constant <= "0000000000000001";
    type_cast_2835_wire_constant <= "0000000000000001";
    type_cast_2860_wire_constant <= "0000000000000000";
    phi_stmt_2649: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2653_wire_constant & type_cast_2655_wire;
      req <= phi_stmt_2649_req_0 & phi_stmt_2649_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2649",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2649_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2649,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2649
    phi_stmt_2656: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2659_wire & type_cast_2661_wire;
      req <= phi_stmt_2656_req_0 & phi_stmt_2656_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2656",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2656_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2656,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2656
    phi_stmt_2715: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2719_wire_constant & type_cast_2721_wire;
      req <= phi_stmt_2715_req_0 & phi_stmt_2715_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2715",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2715_ack_0,
          idata => idata,
          odata => indvar_2715,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2715
    -- flow-through select operator MUX_2862_inst
    input_dim1x_x2_2863 <= type_cast_2860_wire_constant when (cmp88_2847(0) /=  '0') else inc_2837;
    addr_of_2763_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2763_final_reg_req_0;
      addr_of_2763_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2763_final_reg_req_1;
      addr_of_2763_final_reg_ack_1<= rack(0);
      addr_of_2763_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2763_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2762_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_2764,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2793_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2793_final_reg_req_0;
      addr_of_2793_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2793_final_reg_req_1;
      addr_of_2793_final_reg_ack_1<= rack(0);
      addr_of_2793_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2793_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2792_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx70_2794,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2609_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2609_inst_req_0;
      type_cast_2609_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2609_inst_req_1;
      type_cast_2609_inst_ack_1<= rack(0);
      type_cast_2609_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2609_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp12_2523,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv76_2610,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2613_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2613_inst_req_0;
      type_cast_2613_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2613_inst_req_1;
      type_cast_2613_inst_ack_1<= rack(0);
      type_cast_2613_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2613_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp16_2535,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv86_2614,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2623_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2623_inst_req_0;
      type_cast_2623_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2623_inst_req_1;
      type_cast_2623_inst_ack_1<= rack(0);
      type_cast_2623_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2623_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_2505,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv96_2624,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2655_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2655_inst_req_0;
      type_cast_2655_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2655_inst_req_1;
      type_cast_2655_inst_ack_1<= rack(0);
      type_cast_2655_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2655_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2863,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2655_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2659_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2659_inst_req_0;
      type_cast_2659_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2659_inst_req_1;
      type_cast_2659_inst_ack_1<= rack(0);
      type_cast_2659_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2659_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2511,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2659_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2661_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2661_inst_req_0;
      type_cast_2661_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2661_inst_req_1;
      type_cast_2661_inst_ack_1<= rack(0);
      type_cast_2661_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2661_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc92x_xinput_dim0x_x2_2856,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2661_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2721_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2721_inst_req_0;
      type_cast_2721_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2721_inst_req_1;
      type_cast_2721_inst_ack_1<= rack(0);
      type_cast_2721_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2721_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2829,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2721_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2742_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2742_inst_req_0;
      type_cast_2742_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2742_inst_req_1;
      type_cast_2742_inst_ack_1<= rack(0);
      type_cast_2742_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2742_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2741_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv64_2743,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2746_inst
    process(conv64_2743) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv64_2743(31 downto 0);
      type_cast_2746_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2751_inst
    process(ASHR_i32_i32_2750_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2750_wire(31 downto 0);
      shr_2752 <= tmp_var; -- 
    end process;
    type_cast_2756_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2756_inst_req_0;
      type_cast_2756_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2756_inst_req_1;
      type_cast_2756_inst_ack_1<= rack(0);
      type_cast_2756_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2756_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2755_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2757,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2772_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2772_inst_req_0;
      type_cast_2772_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2772_inst_req_1;
      type_cast_2772_inst_ack_1<= rack(0);
      type_cast_2772_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2772_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2771_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv67_2773,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2776_inst
    process(conv67_2773) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv67_2773(31 downto 0);
      type_cast_2776_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2781_inst
    process(ASHR_i32_i32_2780_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2780_wire(31 downto 0);
      shr68_2782 <= tmp_var; -- 
    end process;
    type_cast_2786_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2786_inst_req_0;
      type_cast_2786_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2786_inst_req_1;
      type_cast_2786_inst_ack_1<= rack(0);
      type_cast_2786_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2786_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2785_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom69_2787,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2802_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2802_inst_req_0;
      type_cast_2802_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2802_inst_req_1;
      type_cast_2802_inst_ack_1<= rack(0);
      type_cast_2802_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2802_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2801_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2803,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2812_inst
    process(add74_2809) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add74_2809(31 downto 0);
      type_cast_2812_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2814_inst
    process(conv76_2610) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv76_2610(31 downto 0);
      type_cast_2814_wire <= tmp_var; -- 
    end process;
    type_cast_2841_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2841_inst_req_0;
      type_cast_2841_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2841_inst_req_1;
      type_cast_2841_inst_ack_1<= rack(0);
      type_cast_2841_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2841_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2840_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_2842,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2850_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2850_inst_req_0;
      type_cast_2850_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2850_inst_req_1;
      type_cast_2850_inst_ack_1<= rack(0);
      type_cast_2850_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2850_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp88_2847,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc92_2851,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2867_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2867_inst_req_0;
      type_cast_2867_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2867_inst_req_1;
      type_cast_2867_inst_ack_1<= rack(0);
      type_cast_2867_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2867_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2866_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_2868,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_2559_gather_scatter
    process(LOAD_padding_2559_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_2559_data_0;
      ov(15 downto 0) := iv;
      tmp31_2560 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2762_index_1_rename
    process(R_idxprom_2761_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2761_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2761_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2762_index_1_resize
    process(idxprom_2757) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2757;
      ov := iv(13 downto 0);
      R_idxprom_2761_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2762_root_address_inst
    process(array_obj_ref_2762_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2762_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2762_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2792_index_1_rename
    process(R_idxprom69_2791_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom69_2791_resized;
      ov(13 downto 0) := iv;
      R_idxprom69_2791_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2792_index_1_resize
    process(idxprom69_2787) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom69_2787;
      ov := iv(13 downto 0);
      R_idxprom69_2791_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2792_root_address_inst
    process(array_obj_ref_2792_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2792_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2792_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2504_addr_0
    process(ptr_deref_2504_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2504_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2504_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2504_base_resize
    process(iNsTr_2_2501) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_2501;
      ov := iv(6 downto 0);
      ptr_deref_2504_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2504_gather_scatter
    process(ptr_deref_2504_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2504_data_0;
      ov(15 downto 0) := iv;
      tmp_2505 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2504_root_address_inst
    process(ptr_deref_2504_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2504_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2504_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2522_addr_0
    process(ptr_deref_2522_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2522_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2522_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2522_base_resize
    process(iNsTr_3_2519) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_2519;
      ov := iv(6 downto 0);
      ptr_deref_2522_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2522_gather_scatter
    process(ptr_deref_2522_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2522_data_0;
      ov(15 downto 0) := iv;
      tmp12_2523 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2522_root_address_inst
    process(ptr_deref_2522_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2522_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2522_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2534_addr_0
    process(ptr_deref_2534_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2534_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2534_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2534_base_resize
    process(iNsTr_4_2531) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_2531;
      ov := iv(6 downto 0);
      ptr_deref_2534_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2534_gather_scatter
    process(ptr_deref_2534_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2534_data_0;
      ov(15 downto 0) := iv;
      tmp16_2535 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2534_root_address_inst
    process(ptr_deref_2534_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2534_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2534_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2544_addr_0
    process(ptr_deref_2544_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2544_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2544_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2544_base_resize
    process(iNsTr_5_2541) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_2541;
      ov := iv(0 downto 0);
      ptr_deref_2544_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2544_gather_scatter
    process(ptr_deref_2544_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2544_data_0;
      ov(15 downto 0) := iv;
      tmp25_2545 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2544_root_address_inst
    process(ptr_deref_2544_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2544_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2544_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2556_addr_0
    process(ptr_deref_2556_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2556_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2556_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2556_base_resize
    process(iNsTr_6_2553) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_2553;
      ov := iv(6 downto 0);
      ptr_deref_2556_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2556_gather_scatter
    process(ptr_deref_2556_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2556_data_0;
      ov(15 downto 0) := iv;
      tmp28_2557 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2556_root_address_inst
    process(ptr_deref_2556_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2556_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2556_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2569_addr_0
    process(ptr_deref_2569_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2569_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2569_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2569_base_resize
    process(iNsTr_7_2566) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_2566;
      ov := iv(0 downto 0);
      ptr_deref_2569_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2569_gather_scatter
    process(ptr_deref_2569_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2569_data_0;
      ov(15 downto 0) := iv;
      tmp37_2570 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2569_root_address_inst
    process(ptr_deref_2569_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2569_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2569_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2581_addr_0
    process(ptr_deref_2581_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2581_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2581_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2581_base_resize
    process(iNsTr_8_2578) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_2578;
      ov := iv(6 downto 0);
      ptr_deref_2581_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2581_gather_scatter
    process(ptr_deref_2581_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2581_data_0;
      ov(15 downto 0) := iv;
      tmp40_2582 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2581_root_address_inst
    process(ptr_deref_2581_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2581_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2581_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2593_addr_0
    process(ptr_deref_2593_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2593_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2593_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2593_base_resize
    process(iNsTr_9_2590) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_2590;
      ov := iv(6 downto 0);
      ptr_deref_2593_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2593_gather_scatter
    process(ptr_deref_2593_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2593_data_0;
      ov(15 downto 0) := iv;
      tmp50_2594 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2593_root_address_inst
    process(ptr_deref_2593_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2593_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2593_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2605_addr_0
    process(ptr_deref_2605_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2605_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2605_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2605_base_resize
    process(iNsTr_10_2602) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_2602;
      ov := iv(6 downto 0);
      ptr_deref_2605_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2605_gather_scatter
    process(ptr_deref_2605_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2605_data_0;
      ov(15 downto 0) := iv;
      tmp54_2606 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2605_root_address_inst
    process(ptr_deref_2605_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2605_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2605_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2767_addr_0
    process(ptr_deref_2767_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2767_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2767_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2767_base_resize
    process(arrayidx_2764) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_2764;
      ov := iv(13 downto 0);
      ptr_deref_2767_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2767_gather_scatter
    process(ptr_deref_2767_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2767_data_0;
      ov(63 downto 0) := iv;
      tmp65_2768 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2767_root_address_inst
    process(ptr_deref_2767_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2767_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2767_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2796_addr_0
    process(ptr_deref_2796_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2796_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2796_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2796_base_resize
    process(arrayidx70_2794) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx70_2794;
      ov := iv(13 downto 0);
      ptr_deref_2796_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2796_gather_scatter
    process(tmp65_2768) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp65_2768;
      ov(63 downto 0) := iv;
      ptr_deref_2796_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2796_root_address_inst
    process(ptr_deref_2796_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2796_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2796_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2817_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2816;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2817_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2817_branch_req_0,
          ack0 => if_stmt_2817_branch_ack_0,
          ack1 => if_stmt_2817_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2874_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp97_2873;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2874_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2874_branch_req_0,
          ack0 => if_stmt_2874_branch_ack_0,
          ack1 => if_stmt_2874_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2629_inst
    process(tmp40_2582) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp40_2582, type_cast_2628_wire_constant, tmp_var);
      tmp3_2630 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2640_inst
    process(tmp28_2557) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp28_2557, type_cast_2639_wire_constant, tmp_var);
      tmp7_2641 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2671_inst
    process(input_dim1x_x1x_xph_2649, tmp125_2667) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2649, tmp125_2667, tmp_var);
      tmp126_2672 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2686_inst
    process(tmp4_2635, tmp5_2682) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp4_2635, tmp5_2682, tmp_var);
      tmp6_2687 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2696_inst
    process(tmp8_2646, tmp9_2692) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp8_2646, tmp9_2692, tmp_var);
      tmp10_2697 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2706_inst
    process(tmp6_2687, tmp11_2702) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp6_2687, tmp11_2702, tmp_var);
      tmp13_2707 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2732_inst
    process(tmp127_2677, input_dim2x_x1_2728) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp127_2677, input_dim2x_x1_2728, tmp_var);
      add21_2733 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2737_inst
    process(tmp14_2712, input_dim2x_x1_2728) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp14_2712, input_dim2x_x1_2728, tmp_var);
      add61_2738 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2828_inst
    process(indvar_2715) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2715, type_cast_2827_wire_constant, tmp_var);
      indvarx_xnext_2829 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2836_inst
    process(input_dim1x_x1x_xph_2649) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2649, type_cast_2835_wire_constant, tmp_var);
      inc_2837 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2855_inst
    process(inc92_2851, input_dim0x_x2x_xph_2656) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc92_2851, input_dim0x_x2x_xph_2656, tmp_var);
      inc92x_xinput_dim0x_x2_2856 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2808_inst
    process(conv73_2803) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv73_2803, type_cast_2807_wire_constant, tmp_var);
      add74_2809 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2750_inst
    process(type_cast_2746_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2746_wire, type_cast_2749_wire_constant, tmp_var);
      ASHR_i32_i32_2750_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2780_inst
    process(type_cast_2776_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2776_wire, type_cast_2779_wire_constant, tmp_var);
      ASHR_i32_i32_2780_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2846_inst
    process(conv84_2842, div87_2620) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv84_2842, div87_2620, tmp_var);
      cmp88_2847 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2872_inst
    process(conv94_2868, conv96_2624) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv94_2868, conv96_2624, tmp_var);
      cmp97_2873 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2510_inst
    process(tmp_2505) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_2505, type_cast_2509_wire_constant, tmp_var);
      div_2511 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2619_inst
    process(conv86_2614) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv86_2614, type_cast_2618_wire_constant, tmp_var);
      div87_2620 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2666_inst
    process(tmp16_2535, input_dim0x_x2x_xph_2656) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp16_2535, input_dim0x_x2x_xph_2656, tmp_var);
      tmp125_2667 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2676_inst
    process(tmp12_2523, tmp126_2672) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp12_2523, tmp126_2672, tmp_var);
      tmp127_2677 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2681_inst
    process(tmp37_2570, input_dim1x_x1x_xph_2649) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp37_2570, input_dim1x_x1x_xph_2649, tmp_var);
      tmp5_2682 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2691_inst
    process(tmp25_2545, input_dim0x_x2x_xph_2656) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp25_2545, input_dim0x_x2x_xph_2656, tmp_var);
      tmp9_2692 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2701_inst
    process(tmp54_2606, tmp10_2697) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp54_2606, tmp10_2697, tmp_var);
      tmp11_2702 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2711_inst
    process(tmp50_2594, tmp13_2707) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp50_2594, tmp13_2707, tmp_var);
      tmp14_2712 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2727_inst
    process(indvar_2715) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2715, type_cast_2726_wire_constant, tmp_var);
      input_dim2x_x1_2728 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2815_inst
    process(type_cast_2812_wire, type_cast_2814_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2812_wire, type_cast_2814_wire, tmp_var);
      cmp_2816 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2634_inst
    process(tmp3_2630, tmp31_2560) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp3_2630, tmp31_2560, tmp_var);
      tmp4_2635 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2645_inst
    process(tmp7_2641, tmp31_2560) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp7_2641, tmp31_2560, tmp_var);
      tmp8_2646 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_2762_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2761_scaled;
      array_obj_ref_2762_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2762_index_offset_req_0;
      array_obj_ref_2762_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2762_index_offset_req_1;
      array_obj_ref_2762_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_2792_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom69_2791_scaled;
      array_obj_ref_2792_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2792_index_offset_req_0;
      array_obj_ref_2792_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2792_index_offset_req_1;
      array_obj_ref_2792_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- unary operator type_cast_2741_inst
    process(add21_2733) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add21_2733, tmp_var);
      type_cast_2741_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2755_inst
    process(shr_2752) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2752, tmp_var);
      type_cast_2755_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2771_inst
    process(add61_2738) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add61_2738, tmp_var);
      type_cast_2771_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2785_inst
    process(shr68_2782) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr68_2782, tmp_var);
      type_cast_2785_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2801_inst
    process(input_dim2x_x1_2728) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_2728, tmp_var);
      type_cast_2801_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2840_inst
    process(inc_2837) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2837, tmp_var);
      type_cast_2840_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2866_inst
    process(inc92x_xinput_dim0x_x2_2856) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc92x_xinput_dim0x_x2_2856, tmp_var);
      type_cast_2866_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_2559_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_2559_load_0_req_0;
      LOAD_padding_2559_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_2559_load_0_req_1;
      LOAD_padding_2559_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_2559_word_address_0;
      LOAD_padding_2559_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_2534_load_0 ptr_deref_2522_load_0 ptr_deref_2504_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_2534_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2522_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2504_load_0_req_0;
      ptr_deref_2534_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2522_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2504_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_2534_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2522_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2504_load_0_req_1;
      ptr_deref_2534_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2522_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2504_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2534_word_address_0 & ptr_deref_2522_word_address_0 & ptr_deref_2504_word_address_0;
      ptr_deref_2534_data_0 <= data_out(47 downto 32);
      ptr_deref_2522_data_0 <= data_out(31 downto 16);
      ptr_deref_2504_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 16,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(15 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_2569_load_0 ptr_deref_2544_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2569_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2544_load_0_req_0;
      ptr_deref_2569_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2544_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2569_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2544_load_0_req_1;
      ptr_deref_2569_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2544_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2569_word_address_0 & ptr_deref_2544_word_address_0;
      ptr_deref_2569_data_0 <= data_out(31 downto 16);
      ptr_deref_2544_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(15 downto 0),
          mtag => memory_space_8_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_2556_load_0 ptr_deref_2581_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2556_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2581_load_0_req_0;
      ptr_deref_2556_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2581_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2556_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2581_load_0_req_1;
      ptr_deref_2556_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2581_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2556_word_address_0 & ptr_deref_2581_word_address_0;
      ptr_deref_2556_data_0 <= data_out(31 downto 16);
      ptr_deref_2581_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(15 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_2605_load_0 ptr_deref_2593_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2605_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2593_load_0_req_0;
      ptr_deref_2605_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2593_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2605_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2593_load_0_req_1;
      ptr_deref_2605_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2593_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2605_word_address_0 & ptr_deref_2593_word_address_0;
      ptr_deref_2605_data_0 <= data_out(31 downto 16);
      ptr_deref_2593_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(15 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_2767_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2767_load_0_req_0;
      ptr_deref_2767_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2767_load_0_req_1;
      ptr_deref_2767_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2767_word_address_0;
      ptr_deref_2767_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(13 downto 0),
          mtag => memory_space_4_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(63 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_2796_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2796_store_0_req_0;
      ptr_deref_2796_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2796_store_0_req_1;
      ptr_deref_2796_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2796_word_address_0;
      data_in <= ptr_deref_2796_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(13 downto 0),
          mdata => memory_space_6_sr_data(63 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_start_2491_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_start_2491_inst_req_0;
      RPIPE_Block2_start_2491_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_start_2491_inst_req_1;
      RPIPE_Block2_start_2491_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_2492 <= data_out(15 downto 0);
      Block2_start_read_0_gI: SplitGuardInterface generic map(name => "Block2_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_start_read_0: InputPortRevised -- 
        generic map ( name => "Block2_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_start_pipe_read_req(0),
          oack => Block2_start_pipe_read_ack(0),
          odata => Block2_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2882_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2882_inst_req_0;
      WPIPE_Block2_done_2882_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2882_inst_req_1;
      WPIPE_Block2_done_2882_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_2492;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_8424_start: Boolean;
  signal convTransposeD_CP_8424_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_2905_load_0_req_0 : boolean;
  signal ptr_deref_2905_load_0_ack_0 : boolean;
  signal ptr_deref_2923_load_0_ack_1 : boolean;
  signal ptr_deref_2941_load_0_req_0 : boolean;
  signal ptr_deref_2951_load_0_req_0 : boolean;
  signal RPIPE_Block3_start_2892_inst_req_1 : boolean;
  signal ptr_deref_2941_load_0_ack_1 : boolean;
  signal ptr_deref_2941_load_0_ack_0 : boolean;
  signal RPIPE_Block3_start_2892_inst_ack_1 : boolean;
  signal ptr_deref_2951_load_0_ack_0 : boolean;
  signal ptr_deref_2923_load_0_req_1 : boolean;
  signal ptr_deref_2905_load_0_req_1 : boolean;
  signal RPIPE_Block3_start_2892_inst_req_0 : boolean;
  signal ptr_deref_2941_load_0_req_1 : boolean;
  signal ptr_deref_2923_load_0_req_0 : boolean;
  signal ptr_deref_2923_load_0_ack_0 : boolean;
  signal ptr_deref_2905_load_0_ack_1 : boolean;
  signal RPIPE_Block3_start_2892_inst_ack_0 : boolean;
  signal ptr_deref_2976_load_0_req_0 : boolean;
  signal ptr_deref_2976_load_0_ack_0 : boolean;
  signal ptr_deref_2976_load_0_req_1 : boolean;
  signal ptr_deref_2976_load_0_ack_1 : boolean;
  signal ptr_deref_2963_load_0_req_0 : boolean;
  signal ptr_deref_2963_load_0_ack_0 : boolean;
  signal ptr_deref_2963_load_0_req_1 : boolean;
  signal ptr_deref_2963_load_0_ack_1 : boolean;
  signal ptr_deref_2951_load_0_req_1 : boolean;
  signal ptr_deref_2951_load_0_ack_1 : boolean;
  signal LOAD_padding_2966_load_0_req_0 : boolean;
  signal LOAD_padding_2966_load_0_ack_0 : boolean;
  signal LOAD_padding_2966_load_0_req_1 : boolean;
  signal LOAD_padding_2966_load_0_ack_1 : boolean;
  signal ptr_deref_2988_load_0_req_0 : boolean;
  signal ptr_deref_2988_load_0_ack_0 : boolean;
  signal ptr_deref_2988_load_0_req_1 : boolean;
  signal ptr_deref_2988_load_0_ack_1 : boolean;
  signal ptr_deref_3000_load_0_req_0 : boolean;
  signal ptr_deref_3000_load_0_ack_0 : boolean;
  signal ptr_deref_3000_load_0_req_1 : boolean;
  signal ptr_deref_3000_load_0_ack_1 : boolean;
  signal ptr_deref_3012_load_0_req_0 : boolean;
  signal ptr_deref_3012_load_0_ack_0 : boolean;
  signal ptr_deref_3012_load_0_req_1 : boolean;
  signal ptr_deref_3012_load_0_ack_1 : boolean;
  signal type_cast_3016_inst_req_0 : boolean;
  signal type_cast_3016_inst_ack_0 : boolean;
  signal type_cast_3016_inst_req_1 : boolean;
  signal type_cast_3016_inst_ack_1 : boolean;
  signal type_cast_3020_inst_req_0 : boolean;
  signal type_cast_3020_inst_ack_0 : boolean;
  signal type_cast_3020_inst_req_1 : boolean;
  signal type_cast_3020_inst_ack_1 : boolean;
  signal type_cast_3024_inst_req_0 : boolean;
  signal type_cast_3024_inst_ack_0 : boolean;
  signal type_cast_3024_inst_req_1 : boolean;
  signal type_cast_3024_inst_ack_1 : boolean;
  signal type_cast_3142_inst_req_0 : boolean;
  signal type_cast_3142_inst_ack_0 : boolean;
  signal type_cast_3142_inst_req_1 : boolean;
  signal type_cast_3142_inst_ack_1 : boolean;
  signal type_cast_3156_inst_req_0 : boolean;
  signal type_cast_3156_inst_ack_0 : boolean;
  signal type_cast_3156_inst_req_1 : boolean;
  signal type_cast_3156_inst_ack_1 : boolean;
  signal array_obj_ref_3162_index_offset_req_0 : boolean;
  signal array_obj_ref_3162_index_offset_ack_0 : boolean;
  signal array_obj_ref_3162_index_offset_req_1 : boolean;
  signal array_obj_ref_3162_index_offset_ack_1 : boolean;
  signal addr_of_3163_final_reg_req_0 : boolean;
  signal addr_of_3163_final_reg_ack_0 : boolean;
  signal addr_of_3163_final_reg_req_1 : boolean;
  signal addr_of_3163_final_reg_ack_1 : boolean;
  signal ptr_deref_3167_load_0_req_0 : boolean;
  signal ptr_deref_3167_load_0_ack_0 : boolean;
  signal ptr_deref_3167_load_0_req_1 : boolean;
  signal ptr_deref_3167_load_0_ack_1 : boolean;
  signal type_cast_3172_inst_req_0 : boolean;
  signal type_cast_3172_inst_ack_0 : boolean;
  signal type_cast_3172_inst_req_1 : boolean;
  signal type_cast_3172_inst_ack_1 : boolean;
  signal type_cast_3186_inst_req_0 : boolean;
  signal type_cast_3186_inst_ack_0 : boolean;
  signal type_cast_3186_inst_req_1 : boolean;
  signal type_cast_3186_inst_ack_1 : boolean;
  signal array_obj_ref_3192_index_offset_req_0 : boolean;
  signal array_obj_ref_3192_index_offset_ack_0 : boolean;
  signal array_obj_ref_3192_index_offset_req_1 : boolean;
  signal array_obj_ref_3192_index_offset_ack_1 : boolean;
  signal addr_of_3193_final_reg_req_0 : boolean;
  signal addr_of_3193_final_reg_ack_0 : boolean;
  signal addr_of_3193_final_reg_req_1 : boolean;
  signal addr_of_3193_final_reg_ack_1 : boolean;
  signal ptr_deref_3196_store_0_req_0 : boolean;
  signal ptr_deref_3196_store_0_ack_0 : boolean;
  signal ptr_deref_3196_store_0_req_1 : boolean;
  signal ptr_deref_3196_store_0_ack_1 : boolean;
  signal type_cast_3202_inst_req_0 : boolean;
  signal type_cast_3202_inst_ack_0 : boolean;
  signal type_cast_3202_inst_req_1 : boolean;
  signal type_cast_3202_inst_ack_1 : boolean;
  signal if_stmt_3217_branch_req_0 : boolean;
  signal if_stmt_3217_branch_ack_1 : boolean;
  signal if_stmt_3217_branch_ack_0 : boolean;
  signal type_cast_3241_inst_req_0 : boolean;
  signal type_cast_3241_inst_ack_0 : boolean;
  signal type_cast_3241_inst_req_1 : boolean;
  signal type_cast_3241_inst_ack_1 : boolean;
  signal type_cast_3275_inst_req_0 : boolean;
  signal type_cast_3275_inst_ack_0 : boolean;
  signal type_cast_3275_inst_req_1 : boolean;
  signal type_cast_3275_inst_ack_1 : boolean;
  signal if_stmt_3282_branch_req_0 : boolean;
  signal if_stmt_3282_branch_ack_1 : boolean;
  signal if_stmt_3282_branch_ack_0 : boolean;
  signal WPIPE_Block3_done_3290_inst_req_0 : boolean;
  signal WPIPE_Block3_done_3290_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_3290_inst_req_1 : boolean;
  signal WPIPE_Block3_done_3290_inst_ack_1 : boolean;
  signal type_cast_3053_inst_req_0 : boolean;
  signal type_cast_3053_inst_ack_0 : boolean;
  signal type_cast_3053_inst_req_1 : boolean;
  signal type_cast_3053_inst_ack_1 : boolean;
  signal phi_stmt_3050_req_0 : boolean;
  signal type_cast_3059_inst_req_0 : boolean;
  signal type_cast_3059_inst_ack_0 : boolean;
  signal type_cast_3059_inst_req_1 : boolean;
  signal type_cast_3059_inst_ack_1 : boolean;
  signal phi_stmt_3056_req_0 : boolean;
  signal type_cast_3055_inst_req_0 : boolean;
  signal type_cast_3055_inst_ack_0 : boolean;
  signal type_cast_3055_inst_req_1 : boolean;
  signal type_cast_3055_inst_ack_1 : boolean;
  signal phi_stmt_3050_req_1 : boolean;
  signal type_cast_3061_inst_req_0 : boolean;
  signal type_cast_3061_inst_ack_0 : boolean;
  signal type_cast_3061_inst_req_1 : boolean;
  signal type_cast_3061_inst_ack_1 : boolean;
  signal phi_stmt_3056_req_1 : boolean;
  signal phi_stmt_3050_ack_0 : boolean;
  signal phi_stmt_3056_ack_0 : boolean;
  signal type_cast_3121_inst_req_0 : boolean;
  signal type_cast_3121_inst_ack_0 : boolean;
  signal type_cast_3121_inst_req_1 : boolean;
  signal type_cast_3121_inst_ack_1 : boolean;
  signal phi_stmt_3115_req_1 : boolean;
  signal phi_stmt_3115_req_0 : boolean;
  signal phi_stmt_3115_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_8424_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_8424_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_8424_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_8424_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_8424: Block -- control-path 
    signal convTransposeD_CP_8424_elements: BooleanArray(87 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_8424_elements(0) <= convTransposeD_CP_8424_start;
    convTransposeD_CP_8424_symbol <= convTransposeD_CP_8424_elements(63);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_2890/$entry
      -- CP-element group 0: 	 branch_block_stmt_2890/assign_stmt_2893__entry__
      -- CP-element group 0: 	 branch_block_stmt_2890/assign_stmt_2893/RPIPE_Block3_start_2892_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2890/assign_stmt_2893/RPIPE_Block3_start_2892_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2890/assign_stmt_2893/$entry
      -- CP-element group 0: 	 branch_block_stmt_2890/assign_stmt_2893/RPIPE_Block3_start_2892_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_2890/branch_block_stmt_2890__entry__
      -- CP-element group 0: 	 $entry
      -- 
    rr_8472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(0), ack => RPIPE_Block3_start_2892_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2890/assign_stmt_2893/RPIPE_Block3_start_2892_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_2890/assign_stmt_2893/RPIPE_Block3_start_2892_update_start_
      -- CP-element group 1: 	 branch_block_stmt_2890/assign_stmt_2893/RPIPE_Block3_start_2892_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2890/assign_stmt_2893/RPIPE_Block3_start_2892_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_2890/assign_stmt_2893/RPIPE_Block3_start_2892_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_2890/assign_stmt_2893/RPIPE_Block3_start_2892_Update/$entry
      -- 
    ra_8473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2892_inst_ack_0, ack => convTransposeD_CP_8424_elements(1)); -- 
    cr_8477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(1), ack => RPIPE_Block3_start_2892_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	21 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	6 
    -- CP-element group 2:  members (262) 
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2893__exit__
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2893/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2893/RPIPE_Block3_start_2892_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2893/RPIPE_Block3_start_2892_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2893/RPIPE_Block3_start_2892_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047__entry__
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3016_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3016_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3016_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3020_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3020_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3020_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3024_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3024_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3024_Update/cr
      -- 
    ca_8478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2892_inst_ack_1, ack => convTransposeD_CP_8424_elements(2)); -- 
    rr_8514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => ptr_deref_2905_load_0_req_0); -- 
    rr_8614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => ptr_deref_2941_load_0_req_0); -- 
    rr_8664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => ptr_deref_2951_load_0_req_0); -- 
    cr_8575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => ptr_deref_2923_load_0_req_1); -- 
    cr_8525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => ptr_deref_2905_load_0_req_1); -- 
    cr_8625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => ptr_deref_2941_load_0_req_1); -- 
    rr_8564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => ptr_deref_2923_load_0_req_0); -- 
    rr_8797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => ptr_deref_2976_load_0_req_0); -- 
    cr_8808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => ptr_deref_2976_load_0_req_1); -- 
    rr_8714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => ptr_deref_2963_load_0_req_0); -- 
    cr_8725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => ptr_deref_2963_load_0_req_1); -- 
    cr_8675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => ptr_deref_2951_load_0_req_1); -- 
    rr_8747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => LOAD_padding_2966_load_0_req_0); -- 
    cr_8758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => LOAD_padding_2966_load_0_req_1); -- 
    rr_8847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => ptr_deref_2988_load_0_req_0); -- 
    cr_8858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => ptr_deref_2988_load_0_req_1); -- 
    rr_8897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => ptr_deref_3000_load_0_req_0); -- 
    cr_8908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => ptr_deref_3000_load_0_req_1); -- 
    rr_8947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => ptr_deref_3012_load_0_req_0); -- 
    cr_8958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => ptr_deref_3012_load_0_req_1); -- 
    cr_8977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => type_cast_3016_inst_req_1); -- 
    cr_8991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => type_cast_3020_inst_req_1); -- 
    cr_9005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(2), ack => type_cast_3024_inst_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_Sample/word_access_start/word_0/ra
      -- CP-element group 3: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_Sample/word_access_start/word_0/$exit
      -- 
    ra_8515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2905_load_0_ack_0, ack => convTransposeD_CP_8424_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	27 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_Update/ptr_deref_2905_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_Update/ptr_deref_2905_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_Update/ptr_deref_2905_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2905_Update/ptr_deref_2905_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3024_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3024_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3024_Sample/rr
      -- 
    ca_8526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2905_load_0_ack_1, ack => convTransposeD_CP_8424_elements(4)); -- 
    rr_9000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(4), ack => type_cast_3024_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_Sample/word_access_start/word_0/ra
      -- CP-element group 5: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_sample_completed_
      -- 
    ra_8565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2923_load_0_ack_0, ack => convTransposeD_CP_8424_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	25 
    -- CP-element group 6:  members (12) 
      -- CP-element group 6: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_Update/ptr_deref_2923_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_Update/ptr_deref_2923_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_Update/ptr_deref_2923_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_Update/ptr_deref_2923_Merge/merge_ack
      -- CP-element group 6: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2923_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3020_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3020_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3020_Sample/rr
      -- 
    ca_8576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2923_load_0_ack_1, ack => convTransposeD_CP_8424_elements(6)); -- 
    rr_8986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(6), ack => type_cast_3020_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_Sample/word_access_start/word_0/ra
      -- 
    ra_8615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2941_load_0_ack_0, ack => convTransposeD_CP_8424_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	23 
    -- CP-element group 8:  members (12) 
      -- CP-element group 8: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_Update/ptr_deref_2941_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_Update/ptr_deref_2941_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_Update/ptr_deref_2941_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2941_Update/ptr_deref_2941_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3016_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3016_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3016_Sample/rr
      -- 
    ca_8626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2941_load_0_ack_1, ack => convTransposeD_CP_8424_elements(8)); -- 
    rr_8972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(8), ack => type_cast_3016_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_Sample/word_access_start/word_0/ra
      -- CP-element group 9: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_Sample/word_access_start/$exit
      -- 
    ra_8665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2951_load_0_ack_0, ack => convTransposeD_CP_8424_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	29 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_Update/ptr_deref_2951_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_Update/ptr_deref_2951_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_Update/ptr_deref_2951_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_Update/ptr_deref_2951_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2951_Update/$exit
      -- 
    ca_8676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2951_load_0_ack_1, ack => convTransposeD_CP_8424_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_Sample/word_access_start/word_0/ra
      -- CP-element group 11: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_sample_completed_
      -- 
    ra_8715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2963_load_0_ack_0, ack => convTransposeD_CP_8424_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	29 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_Update/ptr_deref_2963_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_Update/ptr_deref_2963_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_Update/ptr_deref_2963_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_Update/ptr_deref_2963_Merge/merge_ack
      -- CP-element group 12: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2963_update_completed_
      -- 
    ca_8726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2963_load_0_ack_1, ack => convTransposeD_CP_8424_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_Sample/word_access_start/word_0/ra
      -- 
    ra_8748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2966_load_0_ack_0, ack => convTransposeD_CP_8424_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	29 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_Update/LOAD_padding_2966_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_Update/LOAD_padding_2966_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_Update/LOAD_padding_2966_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/LOAD_padding_2966_Update/LOAD_padding_2966_Merge/merge_ack
      -- 
    ca_8759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2966_load_0_ack_1, ack => convTransposeD_CP_8424_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_Sample/word_access_start/word_0/ra
      -- CP-element group 15: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_Sample/word_access_start/word_0/$exit
      -- 
    ra_8798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2976_load_0_ack_0, ack => convTransposeD_CP_8424_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	29 
    -- CP-element group 16:  members (9) 
      -- CP-element group 16: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_Update/ptr_deref_2976_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_Update/ptr_deref_2976_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_Update/ptr_deref_2976_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_Update/ptr_deref_2976_Merge/merge_ack
      -- CP-element group 16: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2976_update_completed_
      -- 
    ca_8809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2976_load_0_ack_1, ack => convTransposeD_CP_8424_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_Sample/word_access_start/word_0/ra
      -- 
    ra_8848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2988_load_0_ack_0, ack => convTransposeD_CP_8424_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	29 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_Update/ptr_deref_2988_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_Update/ptr_deref_2988_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_Update/ptr_deref_2988_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_2988_Update/ptr_deref_2988_Merge/merge_ack
      -- 
    ca_8859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2988_load_0_ack_1, ack => convTransposeD_CP_8424_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_Sample/word_access_start/word_0/ra
      -- 
    ra_8898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3000_load_0_ack_0, ack => convTransposeD_CP_8424_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	29 
    -- CP-element group 20:  members (9) 
      -- CP-element group 20: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_Update/ptr_deref_3000_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_Update/ptr_deref_3000_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_Update/ptr_deref_3000_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3000_Update/ptr_deref_3000_Merge/merge_ack
      -- 
    ca_8909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3000_load_0_ack_1, ack => convTransposeD_CP_8424_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	2 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_Sample/word_access_start/word_0/ra
      -- 
    ra_8948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3012_load_0_ack_0, ack => convTransposeD_CP_8424_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	29 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_Update/word_access_complete/word_0/ca
      -- CP-element group 22: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_Update/ptr_deref_3012_Merge/$entry
      -- CP-element group 22: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_Update/ptr_deref_3012_Merge/$exit
      -- CP-element group 22: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_Update/ptr_deref_3012_Merge/merge_req
      -- CP-element group 22: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/ptr_deref_3012_Update/ptr_deref_3012_Merge/merge_ack
      -- 
    ca_8959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3012_load_0_ack_1, ack => convTransposeD_CP_8424_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3016_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3016_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3016_Sample/ra
      -- 
    ra_8973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3016_inst_ack_0, ack => convTransposeD_CP_8424_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	29 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3016_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3016_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3016_Update/ca
      -- 
    ca_8978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3016_inst_ack_1, ack => convTransposeD_CP_8424_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	6 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3020_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3020_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3020_Sample/ra
      -- 
    ra_8987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3020_inst_ack_0, ack => convTransposeD_CP_8424_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3020_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3020_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3020_Update/ca
      -- 
    ca_8992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3020_inst_ack_1, ack => convTransposeD_CP_8424_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	4 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3024_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3024_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3024_Sample/ra
      -- 
    ra_9001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3024_inst_ack_0, ack => convTransposeD_CP_8424_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3024_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3024_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/type_cast_3024_Update/ca
      -- 
    ca_9006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3024_inst_ack_1, ack => convTransposeD_CP_8424_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  place  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	10 
    -- CP-element group 29: 	12 
    -- CP-element group 29: 	26 
    -- CP-element group 29: 	22 
    -- CP-element group 29: 	14 
    -- CP-element group 29: 	16 
    -- CP-element group 29: 	18 
    -- CP-element group 29: 	20 
    -- CP-element group 29: 	24 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	64 
    -- CP-element group 29: 	65 
    -- CP-element group 29: 	67 
    -- CP-element group 29: 	68 
    -- CP-element group 29:  members (20) 
      -- CP-element group 29: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047__exit__
      -- CP-element group 29: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter
      -- CP-element group 29: 	 branch_block_stmt_2890/assign_stmt_2902_to_assign_stmt_3047/$exit
      -- CP-element group 29: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 29: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/$entry
      -- CP-element group 29: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3053/$entry
      -- CP-element group 29: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3053/SplitProtocol/$entry
      -- CP-element group 29: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3053/SplitProtocol/Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3053/SplitProtocol/Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3053/SplitProtocol/Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3053/SplitProtocol/Update/cr
      -- CP-element group 29: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/$entry
      -- CP-element group 29: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3059/$entry
      -- CP-element group 29: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3059/SplitProtocol/$entry
      -- CP-element group 29: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3059/SplitProtocol/Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3059/SplitProtocol/Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3059/SplitProtocol/Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3059/SplitProtocol/Update/cr
      -- 
    rr_9382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(29), ack => type_cast_3053_inst_req_0); -- 
    cr_9387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(29), ack => type_cast_3053_inst_req_1); -- 
    rr_9405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(29), ack => type_cast_3059_inst_req_0); -- 
    cr_9410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(29), ack => type_cast_3059_inst_req_1); -- 
    convTransposeD_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeD_CP_8424_elements(10) & convTransposeD_CP_8424_elements(12) & convTransposeD_CP_8424_elements(26) & convTransposeD_CP_8424_elements(22) & convTransposeD_CP_8424_elements(14) & convTransposeD_CP_8424_elements(16) & convTransposeD_CP_8424_elements(18) & convTransposeD_CP_8424_elements(20) & convTransposeD_CP_8424_elements(24) & convTransposeD_CP_8424_elements(28);
      gj_convTransposeD_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8424_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	87 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3142_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3142_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3142_Sample/ra
      -- 
    ra_9021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3142_inst_ack_0, ack => convTransposeD_CP_8424_elements(30)); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	87 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3142_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3142_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3142_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3156_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3156_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3156_Sample/rr
      -- 
    ca_9026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3142_inst_ack_1, ack => convTransposeD_CP_8424_elements(31)); -- 
    rr_9034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(31), ack => type_cast_3156_inst_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3156_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3156_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3156_Sample/ra
      -- 
    ra_9035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3156_inst_ack_0, ack => convTransposeD_CP_8424_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	87 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (16) 
      -- CP-element group 33: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3156_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3156_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3156_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_index_resized_1
      -- CP-element group 33: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_index_scaled_1
      -- CP-element group 33: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_index_computed_1
      -- CP-element group 33: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_index_resize_1/$entry
      -- CP-element group 33: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_index_resize_1/$exit
      -- CP-element group 33: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_index_resize_1/index_resize_req
      -- CP-element group 33: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_index_resize_1/index_resize_ack
      -- CP-element group 33: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_index_scale_1/$entry
      -- CP-element group 33: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_index_scale_1/$exit
      -- CP-element group 33: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_index_scale_1/scale_rename_req
      -- CP-element group 33: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_index_scale_1/scale_rename_ack
      -- CP-element group 33: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_final_index_sum_regn_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_final_index_sum_regn_Sample/req
      -- 
    ca_9040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3156_inst_ack_1, ack => convTransposeD_CP_8424_elements(33)); -- 
    req_9065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(33), ack => array_obj_ref_3162_index_offset_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	53 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_final_index_sum_regn_sample_complete
      -- CP-element group 34: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_final_index_sum_regn_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_final_index_sum_regn_Sample/ack
      -- 
    ack_9066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3162_index_offset_ack_0, ack => convTransposeD_CP_8424_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	87 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (11) 
      -- CP-element group 35: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3163_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_root_address_calculated
      -- CP-element group 35: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_offset_calculated
      -- CP-element group 35: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_final_index_sum_regn_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_final_index_sum_regn_Update/ack
      -- CP-element group 35: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_base_plus_offset/$entry
      -- CP-element group 35: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_base_plus_offset/$exit
      -- CP-element group 35: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_base_plus_offset/sum_rename_req
      -- CP-element group 35: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_base_plus_offset/sum_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3163_request/$entry
      -- CP-element group 35: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3163_request/req
      -- 
    ack_9071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3162_index_offset_ack_1, ack => convTransposeD_CP_8424_elements(35)); -- 
    req_9080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(35), ack => addr_of_3163_final_reg_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3163_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3163_request/$exit
      -- CP-element group 36: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3163_request/ack
      -- 
    ack_9081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3163_final_reg_ack_0, ack => convTransposeD_CP_8424_elements(36)); -- 
    -- CP-element group 37:  join  fork  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	87 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (24) 
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3163_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3163_complete/$exit
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3163_complete/ack
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_base_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_word_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_base_address_resized
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_base_addr_resize/$entry
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_base_addr_resize/$exit
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_base_addr_resize/base_resize_req
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_base_addr_resize/base_resize_ack
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_base_plus_offset/$entry
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_base_plus_offset/$exit
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_base_plus_offset/sum_rename_req
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_word_addrgen/$entry
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_word_addrgen/$exit
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_word_addrgen/root_register_req
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_word_addrgen/root_register_ack
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_Sample/word_access_start/$entry
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_Sample/word_access_start/word_0/$entry
      -- CP-element group 37: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_Sample/word_access_start/word_0/rr
      -- 
    ack_9086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3163_final_reg_ack_1, ack => convTransposeD_CP_8424_elements(37)); -- 
    rr_9119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(37), ack => ptr_deref_3167_load_0_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_Sample/word_access_start/$exit
      -- CP-element group 38: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_Sample/word_access_start/word_0/$exit
      -- CP-element group 38: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_Sample/word_access_start/word_0/ra
      -- 
    ra_9120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3167_load_0_ack_0, ack => convTransposeD_CP_8424_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	87 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	48 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_Update/word_access_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_Update/word_access_complete/word_0/$exit
      -- CP-element group 39: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_Update/word_access_complete/word_0/ca
      -- CP-element group 39: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_Update/ptr_deref_3167_Merge/$entry
      -- CP-element group 39: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_Update/ptr_deref_3167_Merge/$exit
      -- CP-element group 39: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_Update/ptr_deref_3167_Merge/merge_req
      -- CP-element group 39: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_Update/ptr_deref_3167_Merge/merge_ack
      -- 
    ca_9131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3167_load_0_ack_1, ack => convTransposeD_CP_8424_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	87 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3172_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3172_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3172_Sample/ra
      -- 
    ra_9145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3172_inst_ack_0, ack => convTransposeD_CP_8424_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	87 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3172_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3172_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3172_Update/ca
      -- CP-element group 41: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3186_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3186_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3186_Sample/rr
      -- 
    ca_9150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3172_inst_ack_1, ack => convTransposeD_CP_8424_elements(41)); -- 
    rr_9158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(41), ack => type_cast_3186_inst_req_0); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3186_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3186_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3186_Sample/ra
      -- 
    ra_9159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3186_inst_ack_0, ack => convTransposeD_CP_8424_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	87 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (16) 
      -- CP-element group 43: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3186_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3186_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3186_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_index_resized_1
      -- CP-element group 43: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_index_scaled_1
      -- CP-element group 43: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_index_computed_1
      -- CP-element group 43: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_index_resize_1/$entry
      -- CP-element group 43: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_index_resize_1/$exit
      -- CP-element group 43: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_index_resize_1/index_resize_req
      -- CP-element group 43: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_index_resize_1/index_resize_ack
      -- CP-element group 43: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_index_scale_1/$entry
      -- CP-element group 43: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_index_scale_1/$exit
      -- CP-element group 43: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_index_scale_1/scale_rename_req
      -- CP-element group 43: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_index_scale_1/scale_rename_ack
      -- CP-element group 43: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_final_index_sum_regn_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_final_index_sum_regn_Sample/req
      -- 
    ca_9164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3186_inst_ack_1, ack => convTransposeD_CP_8424_elements(43)); -- 
    req_9189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(43), ack => array_obj_ref_3192_index_offset_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	53 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_final_index_sum_regn_sample_complete
      -- CP-element group 44: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_final_index_sum_regn_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_final_index_sum_regn_Sample/ack
      -- 
    ack_9190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3192_index_offset_ack_0, ack => convTransposeD_CP_8424_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	87 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (11) 
      -- CP-element group 45: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3193_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_root_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_offset_calculated
      -- CP-element group 45: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_final_index_sum_regn_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_final_index_sum_regn_Update/ack
      -- CP-element group 45: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_base_plus_offset/$entry
      -- CP-element group 45: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_base_plus_offset/$exit
      -- CP-element group 45: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_base_plus_offset/sum_rename_req
      -- CP-element group 45: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_base_plus_offset/sum_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3193_request/$entry
      -- CP-element group 45: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3193_request/req
      -- 
    ack_9195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3192_index_offset_ack_1, ack => convTransposeD_CP_8424_elements(45)); -- 
    req_9204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(45), ack => addr_of_3193_final_reg_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3193_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3193_request/$exit
      -- CP-element group 46: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3193_request/ack
      -- 
    ack_9205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3193_final_reg_ack_0, ack => convTransposeD_CP_8424_elements(46)); -- 
    -- CP-element group 47:  fork  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	87 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (19) 
      -- CP-element group 47: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3193_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3193_complete/$exit
      -- CP-element group 47: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3193_complete/ack
      -- CP-element group 47: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_base_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_word_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_root_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_base_address_resized
      -- CP-element group 47: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_base_addr_resize/$entry
      -- CP-element group 47: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_base_addr_resize/$exit
      -- CP-element group 47: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_base_addr_resize/base_resize_req
      -- CP-element group 47: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_base_addr_resize/base_resize_ack
      -- CP-element group 47: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_base_plus_offset/$entry
      -- CP-element group 47: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_base_plus_offset/$exit
      -- CP-element group 47: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_base_plus_offset/sum_rename_req
      -- CP-element group 47: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_base_plus_offset/sum_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_word_addrgen/$entry
      -- CP-element group 47: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_word_addrgen/$exit
      -- CP-element group 47: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_word_addrgen/root_register_req
      -- CP-element group 47: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_word_addrgen/root_register_ack
      -- 
    ack_9210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3193_final_reg_ack_1, ack => convTransposeD_CP_8424_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	39 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (9) 
      -- CP-element group 48: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_Sample/ptr_deref_3196_Split/$entry
      -- CP-element group 48: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_Sample/ptr_deref_3196_Split/$exit
      -- CP-element group 48: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_Sample/ptr_deref_3196_Split/split_req
      -- CP-element group 48: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_Sample/ptr_deref_3196_Split/split_ack
      -- CP-element group 48: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_Sample/word_access_start/$entry
      -- CP-element group 48: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_Sample/word_access_start/word_0/$entry
      -- CP-element group 48: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_Sample/word_access_start/word_0/rr
      -- 
    rr_9248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(48), ack => ptr_deref_3196_store_0_req_0); -- 
    convTransposeD_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_8424_elements(39) & convTransposeD_CP_8424_elements(47);
      gj_convTransposeD_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8424_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_Sample/word_access_start/$exit
      -- CP-element group 49: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_Sample/word_access_start/word_0/$exit
      -- CP-element group 49: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_Sample/word_access_start/word_0/ra
      -- 
    ra_9249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3196_store_0_ack_0, ack => convTransposeD_CP_8424_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	87 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_Update/word_access_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_Update/word_access_complete/word_0/$exit
      -- CP-element group 50: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_Update/word_access_complete/word_0/ca
      -- 
    ca_9260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3196_store_0_ack_1, ack => convTransposeD_CP_8424_elements(50)); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	87 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3202_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3202_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3202_Sample/ra
      -- 
    ra_9269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3202_inst_ack_0, ack => convTransposeD_CP_8424_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	87 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3202_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3202_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3202_Update/ca
      -- 
    ca_9274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3202_inst_ack_1, ack => convTransposeD_CP_8424_elements(52)); -- 
    -- CP-element group 53:  branch  join  transition  place  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	34 
    -- CP-element group 53: 	52 
    -- CP-element group 53: 	50 
    -- CP-element group 53: 	44 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (10) 
      -- CP-element group 53: 	 branch_block_stmt_2890/if_stmt_3217__entry__
      -- CP-element group 53: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216__exit__
      -- CP-element group 53: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/$exit
      -- CP-element group 53: 	 branch_block_stmt_2890/if_stmt_3217_dead_link/$entry
      -- CP-element group 53: 	 branch_block_stmt_2890/if_stmt_3217_eval_test/$entry
      -- CP-element group 53: 	 branch_block_stmt_2890/if_stmt_3217_eval_test/$exit
      -- CP-element group 53: 	 branch_block_stmt_2890/if_stmt_3217_eval_test/branch_req
      -- CP-element group 53: 	 branch_block_stmt_2890/R_cmp_3218_place
      -- CP-element group 53: 	 branch_block_stmt_2890/if_stmt_3217_if_link/$entry
      -- CP-element group 53: 	 branch_block_stmt_2890/if_stmt_3217_else_link/$entry
      -- 
    branch_req_9282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(53), ack => if_stmt_3217_branch_req_0); -- 
    convTransposeD_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_8424_elements(34) & convTransposeD_CP_8424_elements(52) & convTransposeD_CP_8424_elements(50) & convTransposeD_CP_8424_elements(44);
      gj_convTransposeD_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8424_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	82 
    -- CP-element group 54: 	83 
    -- CP-element group 54:  members (24) 
      -- CP-element group 54: 	 branch_block_stmt_2890/assign_stmt_3229__exit__
      -- CP-element group 54: 	 branch_block_stmt_2890/ifx_xthen_whilex_xbody
      -- CP-element group 54: 	 branch_block_stmt_2890/merge_stmt_3223__exit__
      -- CP-element group 54: 	 branch_block_stmt_2890/assign_stmt_3229__entry__
      -- CP-element group 54: 	 branch_block_stmt_2890/if_stmt_3217_if_link/$exit
      -- CP-element group 54: 	 branch_block_stmt_2890/if_stmt_3217_if_link/if_choice_transition
      -- CP-element group 54: 	 branch_block_stmt_2890/whilex_xbody_ifx_xthen
      -- CP-element group 54: 	 branch_block_stmt_2890/assign_stmt_3229/$entry
      -- CP-element group 54: 	 branch_block_stmt_2890/assign_stmt_3229/$exit
      -- CP-element group 54: 	 branch_block_stmt_2890/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_2890/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3115/$entry
      -- CP-element group 54: 	 branch_block_stmt_2890/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3115/phi_stmt_3115_sources/$entry
      -- CP-element group 54: 	 branch_block_stmt_2890/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3115/phi_stmt_3115_sources/type_cast_3121/$entry
      -- CP-element group 54: 	 branch_block_stmt_2890/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3115/phi_stmt_3115_sources/type_cast_3121/SplitProtocol/$entry
      -- CP-element group 54: 	 branch_block_stmt_2890/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3115/phi_stmt_3115_sources/type_cast_3121/SplitProtocol/Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_2890/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3115/phi_stmt_3115_sources/type_cast_3121/SplitProtocol/Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_2890/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3115/phi_stmt_3115_sources/type_cast_3121/SplitProtocol/Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_2890/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3115/phi_stmt_3115_sources/type_cast_3121/SplitProtocol/Update/cr
      -- CP-element group 54: 	 branch_block_stmt_2890/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_2890/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 54: 	 branch_block_stmt_2890/merge_stmt_3223_PhiReqMerge
      -- CP-element group 54: 	 branch_block_stmt_2890/merge_stmt_3223_PhiAck/$entry
      -- CP-element group 54: 	 branch_block_stmt_2890/merge_stmt_3223_PhiAck/$exit
      -- CP-element group 54: 	 branch_block_stmt_2890/merge_stmt_3223_PhiAck/dummy
      -- 
    if_choice_transition_9287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3217_branch_ack_1, ack => convTransposeD_CP_8424_elements(54)); -- 
    rr_9486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(54), ack => type_cast_3121_inst_req_0); -- 
    cr_9491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(54), ack => type_cast_3121_inst_req_1); -- 
    -- CP-element group 55:  fork  transition  place  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	57 
    -- CP-element group 55: 	59 
    -- CP-element group 55:  members (21) 
      -- CP-element group 55: 	 branch_block_stmt_2890/merge_stmt_3231__exit__
      -- CP-element group 55: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281__entry__
      -- CP-element group 55: 	 branch_block_stmt_2890/merge_stmt_3231_PhiAck/dummy
      -- CP-element group 55: 	 branch_block_stmt_2890/merge_stmt_3231_PhiAck/$exit
      -- CP-element group 55: 	 branch_block_stmt_2890/merge_stmt_3231_PhiReqMerge
      -- CP-element group 55: 	 branch_block_stmt_2890/merge_stmt_3231_PhiAck/$entry
      -- CP-element group 55: 	 branch_block_stmt_2890/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 55: 	 branch_block_stmt_2890/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 55: 	 branch_block_stmt_2890/if_stmt_3217_else_link/$exit
      -- CP-element group 55: 	 branch_block_stmt_2890/if_stmt_3217_else_link/else_choice_transition
      -- CP-element group 55: 	 branch_block_stmt_2890/whilex_xbody_ifx_xelse
      -- CP-element group 55: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/$entry
      -- CP-element group 55: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3241_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3241_update_start_
      -- CP-element group 55: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3241_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3241_Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3241_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3241_Update/cr
      -- CP-element group 55: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3275_update_start_
      -- CP-element group 55: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3275_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3275_Update/cr
      -- 
    else_choice_transition_9291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3217_branch_ack_0, ack => convTransposeD_CP_8424_elements(55)); -- 
    rr_9307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(55), ack => type_cast_3241_inst_req_0); -- 
    cr_9312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(55), ack => type_cast_3241_inst_req_1); -- 
    cr_9326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(55), ack => type_cast_3275_inst_req_1); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3241_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3241_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3241_Sample/ra
      -- 
    ra_9308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3241_inst_ack_0, ack => convTransposeD_CP_8424_elements(56)); -- 
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3241_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3241_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3241_Update/ca
      -- CP-element group 57: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3275_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3275_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3275_Sample/rr
      -- 
    ca_9313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3241_inst_ack_1, ack => convTransposeD_CP_8424_elements(57)); -- 
    rr_9321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(57), ack => type_cast_3275_inst_req_0); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3275_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3275_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3275_Sample/ra
      -- 
    ra_9322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3275_inst_ack_0, ack => convTransposeD_CP_8424_elements(58)); -- 
    -- CP-element group 59:  branch  transition  place  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	55 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (13) 
      -- CP-element group 59: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281__exit__
      -- CP-element group 59: 	 branch_block_stmt_2890/if_stmt_3282__entry__
      -- CP-element group 59: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/$exit
      -- CP-element group 59: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3275_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3275_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_2890/assign_stmt_3237_to_assign_stmt_3281/type_cast_3275_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_2890/if_stmt_3282_dead_link/$entry
      -- CP-element group 59: 	 branch_block_stmt_2890/if_stmt_3282_eval_test/$entry
      -- CP-element group 59: 	 branch_block_stmt_2890/if_stmt_3282_eval_test/$exit
      -- CP-element group 59: 	 branch_block_stmt_2890/if_stmt_3282_eval_test/branch_req
      -- CP-element group 59: 	 branch_block_stmt_2890/R_cmp104_3283_place
      -- CP-element group 59: 	 branch_block_stmt_2890/if_stmt_3282_if_link/$entry
      -- CP-element group 59: 	 branch_block_stmt_2890/if_stmt_3282_else_link/$entry
      -- 
    ca_9327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3275_inst_ack_1, ack => convTransposeD_CP_8424_elements(59)); -- 
    branch_req_9335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(59), ack => if_stmt_3282_branch_req_0); -- 
    -- CP-element group 60:  merge  transition  place  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (15) 
      -- CP-element group 60: 	 branch_block_stmt_2890/merge_stmt_3288__exit__
      -- CP-element group 60: 	 branch_block_stmt_2890/assign_stmt_3292__entry__
      -- CP-element group 60: 	 branch_block_stmt_2890/merge_stmt_3288_PhiReqMerge
      -- CP-element group 60: 	 branch_block_stmt_2890/merge_stmt_3288_PhiAck/dummy
      -- CP-element group 60: 	 branch_block_stmt_2890/merge_stmt_3288_PhiAck/$exit
      -- CP-element group 60: 	 branch_block_stmt_2890/merge_stmt_3288_PhiAck/$entry
      -- CP-element group 60: 	 branch_block_stmt_2890/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_2890/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_2890/if_stmt_3282_if_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_2890/if_stmt_3282_if_link/if_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_2890/ifx_xelse_whilex_xend
      -- CP-element group 60: 	 branch_block_stmt_2890/assign_stmt_3292/$entry
      -- CP-element group 60: 	 branch_block_stmt_2890/assign_stmt_3292/WPIPE_Block3_done_3290_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2890/assign_stmt_3292/WPIPE_Block3_done_3290_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_2890/assign_stmt_3292/WPIPE_Block3_done_3290_Sample/req
      -- 
    if_choice_transition_9340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3282_branch_ack_1, ack => convTransposeD_CP_8424_elements(60)); -- 
    req_9357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(60), ack => WPIPE_Block3_done_3290_inst_req_0); -- 
    -- CP-element group 61:  fork  transition  place  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	71 
    -- CP-element group 61: 	72 
    -- CP-element group 61: 	74 
    -- CP-element group 61: 	75 
    -- CP-element group 61:  members (20) 
      -- CP-element group 61: 	 branch_block_stmt_2890/if_stmt_3282_else_link/$exit
      -- CP-element group 61: 	 branch_block_stmt_2890/if_stmt_3282_else_link/else_choice_transition
      -- CP-element group 61: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 61: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/$entry
      -- CP-element group 61: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3055/$entry
      -- CP-element group 61: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3055/SplitProtocol/$entry
      -- CP-element group 61: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3055/SplitProtocol/Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3055/SplitProtocol/Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3055/SplitProtocol/Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3055/SplitProtocol/Update/cr
      -- CP-element group 61: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/$entry
      -- CP-element group 61: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3061/$entry
      -- CP-element group 61: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3061/SplitProtocol/$entry
      -- CP-element group 61: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3061/SplitProtocol/Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3061/SplitProtocol/Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3061/SplitProtocol/Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3061/SplitProtocol/Update/cr
      -- 
    else_choice_transition_9344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3282_branch_ack_0, ack => convTransposeD_CP_8424_elements(61)); -- 
    rr_9431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(61), ack => type_cast_3055_inst_req_0); -- 
    cr_9436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(61), ack => type_cast_3055_inst_req_1); -- 
    rr_9454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(61), ack => type_cast_3061_inst_req_0); -- 
    cr_9459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(61), ack => type_cast_3061_inst_req_1); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_2890/assign_stmt_3292/WPIPE_Block3_done_3290_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_2890/assign_stmt_3292/WPIPE_Block3_done_3290_update_start_
      -- CP-element group 62: 	 branch_block_stmt_2890/assign_stmt_3292/WPIPE_Block3_done_3290_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_2890/assign_stmt_3292/WPIPE_Block3_done_3290_Sample/ack
      -- CP-element group 62: 	 branch_block_stmt_2890/assign_stmt_3292/WPIPE_Block3_done_3290_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_2890/assign_stmt_3292/WPIPE_Block3_done_3290_Update/req
      -- 
    ack_9358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_3290_inst_ack_0, ack => convTransposeD_CP_8424_elements(62)); -- 
    req_9362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(62), ack => WPIPE_Block3_done_3290_inst_req_1); -- 
    -- CP-element group 63:  transition  place  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (16) 
      -- CP-element group 63: 	 branch_block_stmt_2890/return__
      -- CP-element group 63: 	 branch_block_stmt_2890/assign_stmt_3292__exit__
      -- CP-element group 63: 	 branch_block_stmt_2890/merge_stmt_3294__exit__
      -- CP-element group 63: 	 $exit
      -- CP-element group 63: 	 branch_block_stmt_2890/$exit
      -- CP-element group 63: 	 branch_block_stmt_2890/branch_block_stmt_2890__exit__
      -- CP-element group 63: 	 branch_block_stmt_2890/merge_stmt_3294_PhiAck/dummy
      -- CP-element group 63: 	 branch_block_stmt_2890/merge_stmt_3294_PhiAck/$exit
      -- CP-element group 63: 	 branch_block_stmt_2890/merge_stmt_3294_PhiAck/$entry
      -- CP-element group 63: 	 branch_block_stmt_2890/merge_stmt_3294_PhiReqMerge
      -- CP-element group 63: 	 branch_block_stmt_2890/return___PhiReq/$exit
      -- CP-element group 63: 	 branch_block_stmt_2890/return___PhiReq/$entry
      -- CP-element group 63: 	 branch_block_stmt_2890/assign_stmt_3292/$exit
      -- CP-element group 63: 	 branch_block_stmt_2890/assign_stmt_3292/WPIPE_Block3_done_3290_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_2890/assign_stmt_3292/WPIPE_Block3_done_3290_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_2890/assign_stmt_3292/WPIPE_Block3_done_3290_Update/ack
      -- 
    ack_9363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_3290_inst_ack_1, ack => convTransposeD_CP_8424_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	29 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3053/SplitProtocol/Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3053/SplitProtocol/Sample/ra
      -- 
    ra_9383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3053_inst_ack_0, ack => convTransposeD_CP_8424_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	29 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3053/SplitProtocol/Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3053/SplitProtocol/Update/ca
      -- 
    ca_9388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3053_inst_ack_1, ack => convTransposeD_CP_8424_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	70 
    -- CP-element group 66:  members (5) 
      -- CP-element group 66: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/$exit
      -- CP-element group 66: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/$exit
      -- CP-element group 66: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3053/$exit
      -- CP-element group 66: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3053/SplitProtocol/$exit
      -- CP-element group 66: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_req
      -- 
    phi_stmt_3050_req_9389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3050_req_9389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(66), ack => phi_stmt_3050_req_0); -- 
    convTransposeD_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_8424_elements(64) & convTransposeD_CP_8424_elements(65);
      gj_convTransposeD_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8424_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	29 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3059/SplitProtocol/Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3059/SplitProtocol/Sample/ra
      -- 
    ra_9406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3059_inst_ack_0, ack => convTransposeD_CP_8424_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	29 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3059/SplitProtocol/Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3059/SplitProtocol/Update/ca
      -- 
    ca_9411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3059_inst_ack_1, ack => convTransposeD_CP_8424_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (5) 
      -- CP-element group 69: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/$exit
      -- CP-element group 69: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/$exit
      -- CP-element group 69: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3059/$exit
      -- CP-element group 69: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3059/SplitProtocol/$exit
      -- CP-element group 69: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_req
      -- 
    phi_stmt_3056_req_9412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3056_req_9412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(69), ack => phi_stmt_3056_req_0); -- 
    convTransposeD_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_8424_elements(67) & convTransposeD_CP_8424_elements(68);
      gj_convTransposeD_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8424_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  join  transition  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	66 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	78 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_2890/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_8424_elements(66) & convTransposeD_CP_8424_elements(69);
      gj_convTransposeD_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8424_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	61 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3055/SplitProtocol/Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3055/SplitProtocol/Sample/ra
      -- 
    ra_9432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3055_inst_ack_0, ack => convTransposeD_CP_8424_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	61 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3055/SplitProtocol/Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3055/SplitProtocol/Update/ca
      -- 
    ca_9437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3055_inst_ack_1, ack => convTransposeD_CP_8424_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	77 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/$exit
      -- CP-element group 73: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/$exit
      -- CP-element group 73: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3055/$exit
      -- CP-element group 73: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_sources/type_cast_3055/SplitProtocol/$exit
      -- CP-element group 73: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3050/phi_stmt_3050_req
      -- 
    phi_stmt_3050_req_9438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3050_req_9438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(73), ack => phi_stmt_3050_req_1); -- 
    convTransposeD_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_8424_elements(71) & convTransposeD_CP_8424_elements(72);
      gj_convTransposeD_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8424_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	61 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3061/SplitProtocol/Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3061/SplitProtocol/Sample/ra
      -- 
    ra_9455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3061_inst_ack_0, ack => convTransposeD_CP_8424_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	61 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3061/SplitProtocol/Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3061/SplitProtocol/Update/ca
      -- 
    ca_9460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3061_inst_ack_1, ack => convTransposeD_CP_8424_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/$exit
      -- CP-element group 76: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3061/$exit
      -- CP-element group 76: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_sources/type_cast_3061/SplitProtocol/$exit
      -- CP-element group 76: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_3056/phi_stmt_3056_req
      -- 
    phi_stmt_3056_req_9461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3056_req_9461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(76), ack => phi_stmt_3056_req_1); -- 
    convTransposeD_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_8424_elements(74) & convTransposeD_CP_8424_elements(75);
      gj_convTransposeD_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8424_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	73 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_2890/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_8424_elements(73) & convTransposeD_CP_8424_elements(76);
      gj_convTransposeD_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8424_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  merge  fork  transition  place  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	70 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2890/merge_stmt_3049_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_2890/merge_stmt_3049_PhiAck/$entry
      -- 
    convTransposeD_CP_8424_elements(78) <= OrReduce(convTransposeD_CP_8424_elements(70) & convTransposeD_CP_8424_elements(77));
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_2890/merge_stmt_3049_PhiAck/phi_stmt_3050_ack
      -- 
    phi_stmt_3050_ack_9466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3050_ack_0, ack => convTransposeD_CP_8424_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_2890/merge_stmt_3049_PhiAck/phi_stmt_3056_ack
      -- 
    phi_stmt_3056_ack_9467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3056_ack_0, ack => convTransposeD_CP_8424_elements(80)); -- 
    -- CP-element group 81:  join  transition  place  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (10) 
      -- CP-element group 81: 	 branch_block_stmt_2890/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 81: 	 branch_block_stmt_2890/merge_stmt_3049__exit__
      -- CP-element group 81: 	 branch_block_stmt_2890/assign_stmt_3067_to_assign_stmt_3112__entry__
      -- CP-element group 81: 	 branch_block_stmt_2890/assign_stmt_3067_to_assign_stmt_3112__exit__
      -- CP-element group 81: 	 branch_block_stmt_2890/assign_stmt_3067_to_assign_stmt_3112/$entry
      -- CP-element group 81: 	 branch_block_stmt_2890/assign_stmt_3067_to_assign_stmt_3112/$exit
      -- CP-element group 81: 	 branch_block_stmt_2890/merge_stmt_3049_PhiAck/$exit
      -- CP-element group 81: 	 branch_block_stmt_2890/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 81: 	 branch_block_stmt_2890/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3115/$entry
      -- CP-element group 81: 	 branch_block_stmt_2890/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3115/phi_stmt_3115_sources/$entry
      -- 
    convTransposeD_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_8424_elements(79) & convTransposeD_CP_8424_elements(80);
      gj_convTransposeD_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8424_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	54 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2890/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3115/phi_stmt_3115_sources/type_cast_3121/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2890/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3115/phi_stmt_3115_sources/type_cast_3121/SplitProtocol/Sample/ra
      -- 
    ra_9487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3121_inst_ack_0, ack => convTransposeD_CP_8424_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	54 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2890/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3115/phi_stmt_3115_sources/type_cast_3121/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2890/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3115/phi_stmt_3115_sources/type_cast_3121/SplitProtocol/Update/ca
      -- 
    ca_9492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3121_inst_ack_1, ack => convTransposeD_CP_8424_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (6) 
      -- CP-element group 84: 	 branch_block_stmt_2890/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 84: 	 branch_block_stmt_2890/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3115/$exit
      -- CP-element group 84: 	 branch_block_stmt_2890/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3115/phi_stmt_3115_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2890/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3115/phi_stmt_3115_sources/type_cast_3121/$exit
      -- CP-element group 84: 	 branch_block_stmt_2890/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3115/phi_stmt_3115_sources/type_cast_3121/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2890/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3115/phi_stmt_3115_req
      -- 
    phi_stmt_3115_req_9493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3115_req_9493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(84), ack => phi_stmt_3115_req_1); -- 
    convTransposeD_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_8424_elements(82) & convTransposeD_CP_8424_elements(83);
      gj_convTransposeD_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8424_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  output  delay-element  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	81 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (5) 
      -- CP-element group 85: 	 branch_block_stmt_2890/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 85: 	 branch_block_stmt_2890/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3115/$exit
      -- CP-element group 85: 	 branch_block_stmt_2890/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3115/phi_stmt_3115_sources/$exit
      -- CP-element group 85: 	 branch_block_stmt_2890/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3115/phi_stmt_3115_sources/type_cast_3119_konst_delay_trans
      -- CP-element group 85: 	 branch_block_stmt_2890/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3115/phi_stmt_3115_req
      -- 
    phi_stmt_3115_req_9504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3115_req_9504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(85), ack => phi_stmt_3115_req_0); -- 
    -- Element group convTransposeD_CP_8424_elements(85) is a control-delay.
    cp_element_85_delay: control_delay_element  generic map(name => " 85_delay", delay_value => 1)  port map(req => convTransposeD_CP_8424_elements(81), ack => convTransposeD_CP_8424_elements(85), clk => clk, reset =>reset);
    -- CP-element group 86:  merge  transition  place  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2890/merge_stmt_3114_PhiReqMerge
      -- CP-element group 86: 	 branch_block_stmt_2890/merge_stmt_3114_PhiAck/$entry
      -- 
    convTransposeD_CP_8424_elements(86) <= OrReduce(convTransposeD_CP_8424_elements(85) & convTransposeD_CP_8424_elements(84));
    -- CP-element group 87:  fork  transition  place  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	43 
    -- CP-element group 87: 	35 
    -- CP-element group 87: 	39 
    -- CP-element group 87: 	40 
    -- CP-element group 87: 	41 
    -- CP-element group 87: 	30 
    -- CP-element group 87: 	31 
    -- CP-element group 87: 	33 
    -- CP-element group 87: 	52 
    -- CP-element group 87: 	50 
    -- CP-element group 87: 	51 
    -- CP-element group 87: 	37 
    -- CP-element group 87: 	45 
    -- CP-element group 87: 	47 
    -- CP-element group 87:  members (51) 
      -- CP-element group 87: 	 branch_block_stmt_2890/merge_stmt_3114__exit__
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216__entry__
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/$entry
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3142_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3142_update_start_
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3142_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3142_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3142_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3142_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3156_update_start_
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3156_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3156_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3163_update_start_
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_final_index_sum_regn_update_start
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_final_index_sum_regn_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3162_final_index_sum_regn_Update/req
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3163_complete/$entry
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3163_complete/req
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_update_start_
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_Update/word_access_complete/$entry
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_Update/word_access_complete/word_0/$entry
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3167_Update/word_access_complete/word_0/cr
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3172_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3172_update_start_
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3172_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3172_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3172_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3172_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3186_update_start_
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3186_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3186_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3193_update_start_
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_final_index_sum_regn_update_start
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_final_index_sum_regn_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/array_obj_ref_3192_final_index_sum_regn_Update/req
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3193_complete/$entry
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/addr_of_3193_complete/req
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_update_start_
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_Update/word_access_complete/$entry
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_Update/word_access_complete/word_0/$entry
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/ptr_deref_3196_Update/word_access_complete/word_0/cr
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3202_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3202_update_start_
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3202_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3202_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3202_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_2890/assign_stmt_3128_to_assign_stmt_3216/type_cast_3202_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_2890/merge_stmt_3114_PhiAck/$exit
      -- CP-element group 87: 	 branch_block_stmt_2890/merge_stmt_3114_PhiAck/phi_stmt_3115_ack
      -- 
    phi_stmt_3115_ack_9509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3115_ack_0, ack => convTransposeD_CP_8424_elements(87)); -- 
    rr_9020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(87), ack => type_cast_3142_inst_req_0); -- 
    cr_9025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(87), ack => type_cast_3142_inst_req_1); -- 
    cr_9039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(87), ack => type_cast_3156_inst_req_1); -- 
    req_9070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(87), ack => array_obj_ref_3162_index_offset_req_1); -- 
    req_9085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(87), ack => addr_of_3163_final_reg_req_1); -- 
    cr_9130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(87), ack => ptr_deref_3167_load_0_req_1); -- 
    rr_9144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(87), ack => type_cast_3172_inst_req_0); -- 
    cr_9149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(87), ack => type_cast_3172_inst_req_1); -- 
    cr_9163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(87), ack => type_cast_3186_inst_req_1); -- 
    req_9194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(87), ack => array_obj_ref_3192_index_offset_req_1); -- 
    req_9209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(87), ack => addr_of_3193_final_reg_req_1); -- 
    cr_9259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(87), ack => ptr_deref_3196_store_0_req_1); -- 
    rr_9268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(87), ack => type_cast_3202_inst_req_0); -- 
    cr_9273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8424_elements(87), ack => type_cast_3202_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_3150_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3180_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_2966_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_2966_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom73_3191_resized : std_logic_vector(13 downto 0);
    signal R_idxprom73_3191_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_3161_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_3161_scaled : std_logic_vector(13 downto 0);
    signal add25_3133 : std_logic_vector(15 downto 0);
    signal add65_3138 : std_logic_vector(15 downto 0);
    signal add78_3209 : std_logic_vector(31 downto 0);
    signal array_obj_ref_3162_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3162_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3162_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3162_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3162_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3162_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3192_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3192_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3192_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3192_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3192_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3192_root_address : std_logic_vector(13 downto 0);
    signal arrayidx74_3194 : std_logic_vector(31 downto 0);
    signal arrayidx_3164 : std_logic_vector(31 downto 0);
    signal call_2893 : std_logic_vector(15 downto 0);
    signal cmp104_3281 : std_logic_vector(0 downto 0);
    signal cmp91_3247 : std_logic_vector(0 downto 0);
    signal cmp_3216 : std_logic_vector(0 downto 0);
    signal conv101_3276 : std_logic_vector(31 downto 0);
    signal conv103_3025 : std_logic_vector(31 downto 0);
    signal conv68_3143 : std_logic_vector(31 downto 0);
    signal conv71_3173 : std_logic_vector(31 downto 0);
    signal conv77_3203 : std_logic_vector(31 downto 0);
    signal conv80_3017 : std_logic_vector(31 downto 0);
    signal conv88_3242 : std_logic_vector(31 downto 0);
    signal conv90_3021 : std_logic_vector(31 downto 0);
    signal div5_2930 : std_logic_vector(15 downto 0);
    signal div98_3259 : std_logic_vector(15 downto 0);
    signal div_2912 : std_logic_vector(15 downto 0);
    signal iNsTr_10_3009 : std_logic_vector(31 downto 0);
    signal iNsTr_2_2902 : std_logic_vector(31 downto 0);
    signal iNsTr_3_2920 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2938 : std_logic_vector(31 downto 0);
    signal iNsTr_5_2948 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2960 : std_logic_vector(31 downto 0);
    signal iNsTr_7_2973 : std_logic_vector(31 downto 0);
    signal iNsTr_8_2985 : std_logic_vector(31 downto 0);
    signal iNsTr_9_2997 : std_logic_vector(31 downto 0);
    signal idxprom73_3187 : std_logic_vector(63 downto 0);
    signal idxprom_3157 : std_logic_vector(63 downto 0);
    signal inc95_3253 : std_logic_vector(15 downto 0);
    signal inc_3237 : std_logic_vector(15 downto 0);
    signal indvar_3115 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_3229 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_3271 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_3056 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_3050 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_3265 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_3128 : std_logic_vector(15 downto 0);
    signal ptr_deref_2905_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2905_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2905_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2905_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2905_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2923_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2923_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2923_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2923_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2923_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2941_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2941_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2941_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2941_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2941_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2951_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2951_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2951_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2951_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2951_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2963_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2963_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2963_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2963_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2963_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2976_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2976_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2976_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2976_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2976_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2988_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2988_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2988_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2988_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2988_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3000_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3000_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3000_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3000_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3000_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3012_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3012_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3012_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3012_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3012_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3167_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3167_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3167_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3167_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3167_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3196_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3196_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3196_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3196_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3196_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3196_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr72_3182 : std_logic_vector(31 downto 0);
    signal shr_3152 : std_logic_vector(31 downto 0);
    signal tmp10_3092 : std_logic_vector(15 downto 0);
    signal tmp11_3097 : std_logic_vector(15 downto 0);
    signal tmp12_3102 : std_logic_vector(15 downto 0);
    signal tmp132_3067 : std_logic_vector(15 downto 0);
    signal tmp133_3072 : std_logic_vector(15 downto 0);
    signal tmp134_3077 : std_logic_vector(15 downto 0);
    signal tmp13_3107 : std_logic_vector(15 downto 0);
    signal tmp14_3112 : std_logic_vector(15 downto 0);
    signal tmp16_2942 : std_logic_vector(15 downto 0);
    signal tmp29_2952 : std_logic_vector(15 downto 0);
    signal tmp32_2964 : std_logic_vector(15 downto 0);
    signal tmp35_2967 : std_logic_vector(15 downto 0);
    signal tmp3_2924 : std_logic_vector(15 downto 0);
    signal tmp41_2977 : std_logic_vector(15 downto 0);
    signal tmp44_2989 : std_logic_vector(15 downto 0);
    signal tmp4_3031 : std_logic_vector(15 downto 0);
    signal tmp54_3001 : std_logic_vector(15 downto 0);
    signal tmp58_3013 : std_logic_vector(15 downto 0);
    signal tmp5_3036 : std_logic_vector(15 downto 0);
    signal tmp69_3168 : std_logic_vector(63 downto 0);
    signal tmp6_3082 : std_logic_vector(15 downto 0);
    signal tmp7_3087 : std_logic_vector(15 downto 0);
    signal tmp8_3042 : std_logic_vector(15 downto 0);
    signal tmp9_3047 : std_logic_vector(15 downto 0);
    signal tmp_2906 : std_logic_vector(15 downto 0);
    signal type_cast_2910_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2928_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3029_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3040_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3053_wire : std_logic_vector(15 downto 0);
    signal type_cast_3055_wire : std_logic_vector(15 downto 0);
    signal type_cast_3059_wire : std_logic_vector(15 downto 0);
    signal type_cast_3061_wire : std_logic_vector(15 downto 0);
    signal type_cast_3119_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3121_wire : std_logic_vector(15 downto 0);
    signal type_cast_3126_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3141_wire : std_logic_vector(31 downto 0);
    signal type_cast_3146_wire : std_logic_vector(31 downto 0);
    signal type_cast_3149_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3155_wire : std_logic_vector(63 downto 0);
    signal type_cast_3171_wire : std_logic_vector(31 downto 0);
    signal type_cast_3176_wire : std_logic_vector(31 downto 0);
    signal type_cast_3179_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3185_wire : std_logic_vector(63 downto 0);
    signal type_cast_3201_wire : std_logic_vector(31 downto 0);
    signal type_cast_3207_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3212_wire : std_logic_vector(31 downto 0);
    signal type_cast_3214_wire : std_logic_vector(31 downto 0);
    signal type_cast_3227_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3235_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3240_wire : std_logic_vector(31 downto 0);
    signal type_cast_3251_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3257_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3274_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_2966_word_address_0 <= "0";
    array_obj_ref_3162_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3162_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3162_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3162_resized_base_address <= "00000000000000";
    array_obj_ref_3192_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3192_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3192_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3192_resized_base_address <= "00000000000000";
    iNsTr_10_3009 <= "00000000000000000000000000000101";
    iNsTr_2_2902 <= "00000000000000000000000000000100";
    iNsTr_3_2920 <= "00000000000000000000000000000101";
    iNsTr_4_2938 <= "00000000000000000000000000000110";
    iNsTr_5_2948 <= "00000000000000000000000000000000";
    iNsTr_6_2960 <= "00000000000000000000000000000101";
    iNsTr_7_2973 <= "00000000000000000000000000000001";
    iNsTr_8_2985 <= "00000000000000000000000000000110";
    iNsTr_9_2997 <= "00000000000000000000000000000110";
    ptr_deref_2905_word_offset_0 <= "0000000";
    ptr_deref_2923_word_offset_0 <= "0000000";
    ptr_deref_2941_word_offset_0 <= "0000000";
    ptr_deref_2951_word_offset_0 <= "0";
    ptr_deref_2963_word_offset_0 <= "0000000";
    ptr_deref_2976_word_offset_0 <= "0";
    ptr_deref_2988_word_offset_0 <= "0000000";
    ptr_deref_3000_word_offset_0 <= "0000000";
    ptr_deref_3012_word_offset_0 <= "0000000";
    ptr_deref_3167_word_offset_0 <= "00000000000000";
    ptr_deref_3196_word_offset_0 <= "00000000000000";
    type_cast_2910_wire_constant <= "0000000000000001";
    type_cast_2928_wire_constant <= "0000000000000001";
    type_cast_3029_wire_constant <= "1111111111111111";
    type_cast_3040_wire_constant <= "1111111111111111";
    type_cast_3119_wire_constant <= "0000000000000000";
    type_cast_3126_wire_constant <= "0000000000000100";
    type_cast_3149_wire_constant <= "00000000000000000000000000000010";
    type_cast_3179_wire_constant <= "00000000000000000000000000000010";
    type_cast_3207_wire_constant <= "00000000000000000000000000000100";
    type_cast_3227_wire_constant <= "0000000000000001";
    type_cast_3235_wire_constant <= "0000000000000001";
    type_cast_3251_wire_constant <= "0000000000000001";
    type_cast_3257_wire_constant <= "0000000000000001";
    phi_stmt_3050: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3053_wire & type_cast_3055_wire;
      req <= phi_stmt_3050_req_0 & phi_stmt_3050_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3050",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3050_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_3050,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3050
    phi_stmt_3056: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3059_wire & type_cast_3061_wire;
      req <= phi_stmt_3056_req_0 & phi_stmt_3056_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3056",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3056_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_3056,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3056
    phi_stmt_3115: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3119_wire_constant & type_cast_3121_wire;
      req <= phi_stmt_3115_req_0 & phi_stmt_3115_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3115",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3115_ack_0,
          idata => idata,
          odata => indvar_3115,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3115
    -- flow-through select operator MUX_3264_inst
    input_dim1x_x2_3265 <= div98_3259 when (cmp91_3247(0) /=  '0') else inc_3237;
    -- flow-through select operator MUX_3270_inst
    input_dim0x_x0_3271 <= inc95_3253 when (cmp91_3247(0) /=  '0') else input_dim0x_x2x_xph_3056;
    addr_of_3163_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3163_final_reg_req_0;
      addr_of_3163_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3163_final_reg_req_1;
      addr_of_3163_final_reg_ack_1<= rack(0);
      addr_of_3163_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3163_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3162_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_3164,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3193_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3193_final_reg_req_0;
      addr_of_3193_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3193_final_reg_req_1;
      addr_of_3193_final_reg_ack_1<= rack(0);
      addr_of_3193_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3193_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3192_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx74_3194,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3016_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3016_inst_req_0;
      type_cast_3016_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3016_inst_req_1;
      type_cast_3016_inst_ack_1<= rack(0);
      type_cast_3016_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3016_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp16_2942,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv80_3017,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3020_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3020_inst_req_0;
      type_cast_3020_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3020_inst_req_1;
      type_cast_3020_inst_ack_1<= rack(0);
      type_cast_3020_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3020_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3_2924,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_3021,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3024_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3024_inst_req_0;
      type_cast_3024_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3024_inst_req_1;
      type_cast_3024_inst_ack_1<= rack(0);
      type_cast_3024_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3024_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_2906,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv103_3025,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3053_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3053_inst_req_0;
      type_cast_3053_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3053_inst_req_1;
      type_cast_3053_inst_ack_1<= rack(0);
      type_cast_3053_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3053_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div5_2930,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3053_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3055_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3055_inst_req_0;
      type_cast_3055_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3055_inst_req_1;
      type_cast_3055_inst_ack_1<= rack(0);
      type_cast_3055_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3055_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_3265,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3055_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3059_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3059_inst_req_0;
      type_cast_3059_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3059_inst_req_1;
      type_cast_3059_inst_ack_1<= rack(0);
      type_cast_3059_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3059_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2912,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3059_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3061_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3061_inst_req_0;
      type_cast_3061_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3061_inst_req_1;
      type_cast_3061_inst_ack_1<= rack(0);
      type_cast_3061_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3061_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_3271,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3061_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3121_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3121_inst_req_0;
      type_cast_3121_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3121_inst_req_1;
      type_cast_3121_inst_ack_1<= rack(0);
      type_cast_3121_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3121_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_3229,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3121_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3142_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3142_inst_req_0;
      type_cast_3142_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3142_inst_req_1;
      type_cast_3142_inst_ack_1<= rack(0);
      type_cast_3142_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3142_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3141_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_3143,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3146_inst
    process(conv68_3143) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv68_3143(31 downto 0);
      type_cast_3146_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3151_inst
    process(ASHR_i32_i32_3150_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3150_wire(31 downto 0);
      shr_3152 <= tmp_var; -- 
    end process;
    type_cast_3156_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3156_inst_req_0;
      type_cast_3156_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3156_inst_req_1;
      type_cast_3156_inst_ack_1<= rack(0);
      type_cast_3156_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3156_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3155_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_3157,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3172_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3172_inst_req_0;
      type_cast_3172_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3172_inst_req_1;
      type_cast_3172_inst_ack_1<= rack(0);
      type_cast_3172_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3172_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3171_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_3173,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3176_inst
    process(conv71_3173) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv71_3173(31 downto 0);
      type_cast_3176_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3181_inst
    process(ASHR_i32_i32_3180_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3180_wire(31 downto 0);
      shr72_3182 <= tmp_var; -- 
    end process;
    type_cast_3186_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3186_inst_req_0;
      type_cast_3186_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3186_inst_req_1;
      type_cast_3186_inst_ack_1<= rack(0);
      type_cast_3186_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3186_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3185_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom73_3187,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3202_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3202_inst_req_0;
      type_cast_3202_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3202_inst_req_1;
      type_cast_3202_inst_ack_1<= rack(0);
      type_cast_3202_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3202_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3201_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv77_3203,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3212_inst
    process(add78_3209) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add78_3209(31 downto 0);
      type_cast_3212_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3214_inst
    process(conv80_3017) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv80_3017(31 downto 0);
      type_cast_3214_wire <= tmp_var; -- 
    end process;
    type_cast_3241_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3241_inst_req_0;
      type_cast_3241_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3241_inst_req_1;
      type_cast_3241_inst_ack_1<= rack(0);
      type_cast_3241_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3241_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3240_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv88_3242,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3275_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3275_inst_req_0;
      type_cast_3275_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3275_inst_req_1;
      type_cast_3275_inst_ack_1<= rack(0);
      type_cast_3275_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3275_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3274_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv101_3276,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_2966_gather_scatter
    process(LOAD_padding_2966_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_2966_data_0;
      ov(15 downto 0) := iv;
      tmp35_2967 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3162_index_1_rename
    process(R_idxprom_3161_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_3161_resized;
      ov(13 downto 0) := iv;
      R_idxprom_3161_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3162_index_1_resize
    process(idxprom_3157) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_3157;
      ov := iv(13 downto 0);
      R_idxprom_3161_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3162_root_address_inst
    process(array_obj_ref_3162_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3162_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3162_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3192_index_1_rename
    process(R_idxprom73_3191_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom73_3191_resized;
      ov(13 downto 0) := iv;
      R_idxprom73_3191_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3192_index_1_resize
    process(idxprom73_3187) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom73_3187;
      ov := iv(13 downto 0);
      R_idxprom73_3191_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3192_root_address_inst
    process(array_obj_ref_3192_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3192_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3192_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2905_addr_0
    process(ptr_deref_2905_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2905_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2905_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2905_base_resize
    process(iNsTr_2_2902) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_2902;
      ov := iv(6 downto 0);
      ptr_deref_2905_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2905_gather_scatter
    process(ptr_deref_2905_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2905_data_0;
      ov(15 downto 0) := iv;
      tmp_2906 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2905_root_address_inst
    process(ptr_deref_2905_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2905_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2905_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2923_addr_0
    process(ptr_deref_2923_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2923_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2923_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2923_base_resize
    process(iNsTr_3_2920) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_2920;
      ov := iv(6 downto 0);
      ptr_deref_2923_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2923_gather_scatter
    process(ptr_deref_2923_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2923_data_0;
      ov(15 downto 0) := iv;
      tmp3_2924 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2923_root_address_inst
    process(ptr_deref_2923_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2923_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2923_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2941_addr_0
    process(ptr_deref_2941_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2941_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2941_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2941_base_resize
    process(iNsTr_4_2938) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_2938;
      ov := iv(6 downto 0);
      ptr_deref_2941_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2941_gather_scatter
    process(ptr_deref_2941_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2941_data_0;
      ov(15 downto 0) := iv;
      tmp16_2942 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2941_root_address_inst
    process(ptr_deref_2941_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2941_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2941_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2951_addr_0
    process(ptr_deref_2951_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2951_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2951_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2951_base_resize
    process(iNsTr_5_2948) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_2948;
      ov := iv(0 downto 0);
      ptr_deref_2951_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2951_gather_scatter
    process(ptr_deref_2951_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2951_data_0;
      ov(15 downto 0) := iv;
      tmp29_2952 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2951_root_address_inst
    process(ptr_deref_2951_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2951_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2951_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2963_addr_0
    process(ptr_deref_2963_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2963_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2963_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2963_base_resize
    process(iNsTr_6_2960) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_2960;
      ov := iv(6 downto 0);
      ptr_deref_2963_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2963_gather_scatter
    process(ptr_deref_2963_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2963_data_0;
      ov(15 downto 0) := iv;
      tmp32_2964 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2963_root_address_inst
    process(ptr_deref_2963_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2963_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2963_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2976_addr_0
    process(ptr_deref_2976_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2976_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2976_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2976_base_resize
    process(iNsTr_7_2973) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_2973;
      ov := iv(0 downto 0);
      ptr_deref_2976_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2976_gather_scatter
    process(ptr_deref_2976_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2976_data_0;
      ov(15 downto 0) := iv;
      tmp41_2977 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2976_root_address_inst
    process(ptr_deref_2976_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2976_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2976_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2988_addr_0
    process(ptr_deref_2988_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2988_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2988_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2988_base_resize
    process(iNsTr_8_2985) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_2985;
      ov := iv(6 downto 0);
      ptr_deref_2988_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2988_gather_scatter
    process(ptr_deref_2988_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2988_data_0;
      ov(15 downto 0) := iv;
      tmp44_2989 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2988_root_address_inst
    process(ptr_deref_2988_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2988_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2988_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3000_addr_0
    process(ptr_deref_3000_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3000_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_3000_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3000_base_resize
    process(iNsTr_9_2997) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_2997;
      ov := iv(6 downto 0);
      ptr_deref_3000_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3000_gather_scatter
    process(ptr_deref_3000_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3000_data_0;
      ov(15 downto 0) := iv;
      tmp54_3001 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3000_root_address_inst
    process(ptr_deref_3000_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3000_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_3000_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3012_addr_0
    process(ptr_deref_3012_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3012_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_3012_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3012_base_resize
    process(iNsTr_10_3009) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_3009;
      ov := iv(6 downto 0);
      ptr_deref_3012_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3012_gather_scatter
    process(ptr_deref_3012_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3012_data_0;
      ov(15 downto 0) := iv;
      tmp58_3013 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3012_root_address_inst
    process(ptr_deref_3012_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3012_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_3012_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3167_addr_0
    process(ptr_deref_3167_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3167_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3167_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3167_base_resize
    process(arrayidx_3164) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_3164;
      ov := iv(13 downto 0);
      ptr_deref_3167_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3167_gather_scatter
    process(ptr_deref_3167_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3167_data_0;
      ov(63 downto 0) := iv;
      tmp69_3168 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3167_root_address_inst
    process(ptr_deref_3167_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3167_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3167_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3196_addr_0
    process(ptr_deref_3196_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3196_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3196_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3196_base_resize
    process(arrayidx74_3194) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx74_3194;
      ov := iv(13 downto 0);
      ptr_deref_3196_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3196_gather_scatter
    process(tmp69_3168) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp69_3168;
      ov(63 downto 0) := iv;
      ptr_deref_3196_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3196_root_address_inst
    process(ptr_deref_3196_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3196_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3196_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_3217_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_3216;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3217_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3217_branch_req_0,
          ack0 => if_stmt_3217_branch_ack_0,
          ack1 => if_stmt_3217_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3282_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp104_3281;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3282_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3282_branch_req_0,
          ack0 => if_stmt_3282_branch_ack_0,
          ack1 => if_stmt_3282_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_3030_inst
    process(tmp44_2989) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp44_2989, type_cast_3029_wire_constant, tmp_var);
      tmp4_3031 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3041_inst
    process(tmp32_2964) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp32_2964, type_cast_3040_wire_constant, tmp_var);
      tmp8_3042 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3071_inst
    process(input_dim1x_x1x_xph_3050, tmp132_3067) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_3050, tmp132_3067, tmp_var);
      tmp133_3072 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3086_inst
    process(tmp5_3036, tmp6_3082) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp5_3036, tmp6_3082, tmp_var);
      tmp7_3087 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3096_inst
    process(tmp9_3047, tmp10_3092) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp9_3047, tmp10_3092, tmp_var);
      tmp11_3097 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3106_inst
    process(tmp7_3087, tmp12_3102) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp7_3087, tmp12_3102, tmp_var);
      tmp13_3107 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3132_inst
    process(tmp134_3077, input_dim2x_x1_3128) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp134_3077, input_dim2x_x1_3128, tmp_var);
      add25_3133 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3137_inst
    process(tmp14_3112, input_dim2x_x1_3128) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp14_3112, input_dim2x_x1_3128, tmp_var);
      add65_3138 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3228_inst
    process(indvar_3115) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_3115, type_cast_3227_wire_constant, tmp_var);
      indvarx_xnext_3229 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3236_inst
    process(input_dim1x_x1x_xph_3050) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_3050, type_cast_3235_wire_constant, tmp_var);
      inc_3237 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3252_inst
    process(input_dim0x_x2x_xph_3056) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim0x_x2x_xph_3056, type_cast_3251_wire_constant, tmp_var);
      inc95_3253 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3208_inst
    process(conv77_3203) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv77_3203, type_cast_3207_wire_constant, tmp_var);
      add78_3209 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3150_inst
    process(type_cast_3146_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3146_wire, type_cast_3149_wire_constant, tmp_var);
      ASHR_i32_i32_3150_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3180_inst
    process(type_cast_3176_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3176_wire, type_cast_3179_wire_constant, tmp_var);
      ASHR_i32_i32_3180_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3246_inst
    process(conv88_3242, conv90_3021) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv88_3242, conv90_3021, tmp_var);
      cmp91_3247 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3280_inst
    process(conv101_3276, conv103_3025) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv101_3276, conv103_3025, tmp_var);
      cmp104_3281 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2911_inst
    process(tmp_2906) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_2906, type_cast_2910_wire_constant, tmp_var);
      div_2912 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2929_inst
    process(tmp3_2924) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp3_2924, type_cast_2928_wire_constant, tmp_var);
      div5_2930 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_3258_inst
    process(tmp3_2924) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp3_2924, type_cast_3257_wire_constant, tmp_var);
      div98_3259 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3066_inst
    process(tmp3_2924, input_dim0x_x2x_xph_3056) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp3_2924, input_dim0x_x2x_xph_3056, tmp_var);
      tmp132_3067 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3076_inst
    process(tmp16_2942, tmp133_3072) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp16_2942, tmp133_3072, tmp_var);
      tmp134_3077 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3081_inst
    process(tmp41_2977, input_dim1x_x1x_xph_3050) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp41_2977, input_dim1x_x1x_xph_3050, tmp_var);
      tmp6_3082 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3091_inst
    process(tmp29_2952, input_dim0x_x2x_xph_3056) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp29_2952, input_dim0x_x2x_xph_3056, tmp_var);
      tmp10_3092 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3101_inst
    process(tmp58_3013, tmp11_3097) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp58_3013, tmp11_3097, tmp_var);
      tmp12_3102 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3111_inst
    process(tmp54_3001, tmp13_3107) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp54_3001, tmp13_3107, tmp_var);
      tmp14_3112 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3127_inst
    process(indvar_3115) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_3115, type_cast_3126_wire_constant, tmp_var);
      input_dim2x_x1_3128 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3215_inst
    process(type_cast_3212_wire, type_cast_3214_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3212_wire, type_cast_3214_wire, tmp_var);
      cmp_3216 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_3035_inst
    process(tmp4_3031, tmp35_2967) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp4_3031, tmp35_2967, tmp_var);
      tmp5_3036 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_3046_inst
    process(tmp8_3042, tmp35_2967) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp8_3042, tmp35_2967, tmp_var);
      tmp9_3047 <= tmp_var; --
    end process;
    -- shared split operator group (29) : array_obj_ref_3162_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_3161_scaled;
      array_obj_ref_3162_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3162_index_offset_req_0;
      array_obj_ref_3162_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3162_index_offset_req_1;
      array_obj_ref_3162_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : array_obj_ref_3192_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom73_3191_scaled;
      array_obj_ref_3192_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3192_index_offset_req_0;
      array_obj_ref_3192_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3192_index_offset_req_1;
      array_obj_ref_3192_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- unary operator type_cast_3141_inst
    process(add25_3133) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add25_3133, tmp_var);
      type_cast_3141_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3155_inst
    process(shr_3152) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_3152, tmp_var);
      type_cast_3155_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3171_inst
    process(add65_3138) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add65_3138, tmp_var);
      type_cast_3171_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3185_inst
    process(shr72_3182) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr72_3182, tmp_var);
      type_cast_3185_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3201_inst
    process(input_dim2x_x1_3128) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_3128, tmp_var);
      type_cast_3201_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3240_inst
    process(inc_3237) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_3237, tmp_var);
      type_cast_3240_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3274_inst
    process(input_dim0x_x0_3271) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x0_3271, tmp_var);
      type_cast_3274_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_2966_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_2966_load_0_req_0;
      LOAD_padding_2966_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_2966_load_0_req_1;
      LOAD_padding_2966_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_2966_word_address_0;
      LOAD_padding_2966_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_2941_load_0 ptr_deref_2923_load_0 ptr_deref_2905_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_2941_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2923_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2905_load_0_req_0;
      ptr_deref_2941_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2923_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2905_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_2941_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2923_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2905_load_0_req_1;
      ptr_deref_2941_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2923_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2905_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2941_word_address_0 & ptr_deref_2923_word_address_0 & ptr_deref_2905_word_address_0;
      ptr_deref_2941_data_0 <= data_out(47 downto 32);
      ptr_deref_2923_data_0 <= data_out(31 downto 16);
      ptr_deref_2905_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 16,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(15 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_2976_load_0 ptr_deref_2951_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2976_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2951_load_0_req_0;
      ptr_deref_2976_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2951_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2976_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2951_load_0_req_1;
      ptr_deref_2976_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2951_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2976_word_address_0 & ptr_deref_2951_word_address_0;
      ptr_deref_2976_data_0 <= data_out(31 downto 16);
      ptr_deref_2951_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(15 downto 0),
          mtag => memory_space_8_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_2963_load_0 ptr_deref_2988_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2963_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2988_load_0_req_0;
      ptr_deref_2963_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2988_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2963_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2988_load_0_req_1;
      ptr_deref_2963_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2988_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2963_word_address_0 & ptr_deref_2988_word_address_0;
      ptr_deref_2963_data_0 <= data_out(31 downto 16);
      ptr_deref_2988_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(15 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_3000_load_0 ptr_deref_3012_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_3000_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_3012_load_0_req_0;
      ptr_deref_3000_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_3012_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_3000_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_3012_load_0_req_1;
      ptr_deref_3000_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_3012_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_3000_word_address_0 & ptr_deref_3012_word_address_0;
      ptr_deref_3000_data_0 <= data_out(31 downto 16);
      ptr_deref_3012_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(15 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_3167_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_3167_load_0_req_0;
      ptr_deref_3167_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_3167_load_0_req_1;
      ptr_deref_3167_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_3167_word_address_0;
      ptr_deref_3167_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(13 downto 0),
          mtag => memory_space_4_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(63 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_3196_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_3196_store_0_req_0;
      ptr_deref_3196_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_3196_store_0_req_1;
      ptr_deref_3196_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_3196_word_address_0;
      data_in <= ptr_deref_3196_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(13 downto 0),
          mdata => memory_space_6_sr_data(63 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_start_2892_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_start_2892_inst_req_0;
      RPIPE_Block3_start_2892_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_start_2892_inst_req_1;
      RPIPE_Block3_start_2892_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_2893 <= data_out(15 downto 0);
      Block3_start_read_0_gI: SplitGuardInterface generic map(name => "Block3_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_start_read_0: InputPortRevised -- 
        generic map ( name => "Block3_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_start_pipe_read_req(0),
          oack => Block3_start_pipe_read_ack(0),
          odata => Block3_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_3290_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_3290_inst_req_0;
      WPIPE_Block3_done_3290_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_3290_inst_req_1;
      WPIPE_Block3_done_3290_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_2893;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendOutput is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendOutput;
architecture sendOutput_arch of sendOutput is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal sendOutput_CP_4163_start: Boolean;
  signal sendOutput_CP_4163_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1541_inst_ack_0 : boolean;
  signal array_obj_ref_1492_index_offset_ack_1 : boolean;
  signal array_obj_ref_1492_index_offset_req_1 : boolean;
  signal type_cast_1531_inst_ack_1 : boolean;
  signal if_stmt_1436_branch_ack_1 : boolean;
  signal array_obj_ref_1492_index_offset_ack_0 : boolean;
  signal type_cast_1531_inst_req_1 : boolean;
  signal type_cast_1521_inst_req_1 : boolean;
  signal ptr_deref_1414_load_0_req_0 : boolean;
  signal type_cast_1511_inst_req_1 : boolean;
  signal type_cast_1531_inst_req_0 : boolean;
  signal if_stmt_1436_branch_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1573_inst_req_1 : boolean;
  signal type_cast_1511_inst_req_0 : boolean;
  signal ptr_deref_1497_load_0_ack_0 : boolean;
  signal type_cast_1571_inst_ack_0 : boolean;
  signal type_cast_1501_inst_ack_1 : boolean;
  signal addr_of_1493_final_reg_req_0 : boolean;
  signal array_obj_ref_1492_index_offset_req_0 : boolean;
  signal type_cast_1561_inst_ack_0 : boolean;
  signal type_cast_1501_inst_req_1 : boolean;
  signal type_cast_1511_inst_ack_1 : boolean;
  signal type_cast_1418_inst_ack_0 : boolean;
  signal ptr_deref_1414_load_0_req_1 : boolean;
  signal type_cast_1551_inst_ack_0 : boolean;
  signal type_cast_1418_inst_req_1 : boolean;
  signal type_cast_1402_inst_req_0 : boolean;
  signal type_cast_1561_inst_req_0 : boolean;
  signal type_cast_1571_inst_ack_1 : boolean;
  signal ptr_deref_1497_load_0_req_0 : boolean;
  signal type_cast_1501_inst_ack_0 : boolean;
  signal type_cast_1501_inst_req_0 : boolean;
  signal type_cast_1561_inst_ack_1 : boolean;
  signal type_cast_1402_inst_req_1 : boolean;
  signal type_cast_1571_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1573_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1573_inst_req_0 : boolean;
  signal type_cast_1541_inst_ack_1 : boolean;
  signal type_cast_1402_inst_ack_1 : boolean;
  signal type_cast_1418_inst_ack_1 : boolean;
  signal type_cast_1463_inst_req_0 : boolean;
  signal type_cast_1463_inst_ack_1 : boolean;
  signal type_cast_1551_inst_req_0 : boolean;
  signal type_cast_1521_inst_ack_0 : boolean;
  signal type_cast_1511_inst_ack_0 : boolean;
  signal type_cast_1551_inst_ack_1 : boolean;
  signal type_cast_1551_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1573_inst_ack_0 : boolean;
  signal type_cast_1521_inst_req_0 : boolean;
  signal type_cast_1402_inst_ack_0 : boolean;
  signal type_cast_1531_inst_ack_0 : boolean;
  signal ptr_deref_1414_load_0_ack_0 : boolean;
  signal type_cast_1541_inst_req_1 : boolean;
  signal type_cast_1571_inst_req_0 : boolean;
  signal type_cast_1463_inst_req_1 : boolean;
  signal type_cast_1561_inst_req_1 : boolean;
  signal addr_of_1493_final_reg_ack_0 : boolean;
  signal ptr_deref_1497_load_0_req_1 : boolean;
  signal type_cast_1418_inst_req_0 : boolean;
  signal type_cast_1541_inst_req_0 : boolean;
  signal type_cast_1521_inst_ack_1 : boolean;
  signal ptr_deref_1414_load_0_ack_1 : boolean;
  signal if_stmt_1436_branch_ack_0 : boolean;
  signal ptr_deref_1497_load_0_ack_1 : boolean;
  signal type_cast_1463_inst_ack_0 : boolean;
  signal addr_of_1493_final_reg_ack_1 : boolean;
  signal addr_of_1493_final_reg_req_1 : boolean;
  signal ptr_deref_1382_load_0_req_0 : boolean;
  signal ptr_deref_1382_load_0_ack_0 : boolean;
  signal ptr_deref_1382_load_0_req_1 : boolean;
  signal ptr_deref_1382_load_0_ack_1 : boolean;
  signal type_cast_1386_inst_req_0 : boolean;
  signal type_cast_1386_inst_ack_0 : boolean;
  signal type_cast_1386_inst_req_1 : boolean;
  signal type_cast_1386_inst_ack_1 : boolean;
  signal ptr_deref_1398_load_0_req_0 : boolean;
  signal ptr_deref_1398_load_0_ack_0 : boolean;
  signal ptr_deref_1398_load_0_req_1 : boolean;
  signal ptr_deref_1398_load_0_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1576_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1576_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1576_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1576_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1579_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1579_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1579_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1579_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1582_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1582_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1582_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1582_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1585_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1585_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1585_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1585_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1588_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1588_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1588_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1588_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1591_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1591_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1591_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1591_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1594_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1594_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1594_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1594_inst_ack_1 : boolean;
  signal if_stmt_1608_branch_req_0 : boolean;
  signal if_stmt_1608_branch_ack_1 : boolean;
  signal if_stmt_1608_branch_ack_0 : boolean;
  signal phi_stmt_1480_req_0 : boolean;
  signal type_cast_1486_inst_req_0 : boolean;
  signal type_cast_1486_inst_ack_0 : boolean;
  signal type_cast_1486_inst_req_1 : boolean;
  signal type_cast_1486_inst_ack_1 : boolean;
  signal phi_stmt_1480_req_1 : boolean;
  signal phi_stmt_1480_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendOutput_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendOutput_CP_4163_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendOutput_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_4163_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendOutput_CP_4163_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_4163_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendOutput_CP_4163: Block -- control-path 
    signal sendOutput_CP_4163_elements: BooleanArray(72 downto 0);
    -- 
  begin -- 
    sendOutput_CP_4163_elements(0) <= sendOutput_CP_4163_start;
    sendOutput_CP_4163_symbol <= sendOutput_CP_4163_elements(72);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	10 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	8 
    -- CP-element group 0:  members (92) 
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1418_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1418_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1402_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1418_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1402_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1371/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/branch_block_stmt_1371__entry__
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435__entry__
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1386_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1386_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1386_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1402_update_start_
      -- 
    rr_4354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(0), ack => ptr_deref_1414_load_0_req_0); -- 
    cr_4365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(0), ack => ptr_deref_1414_load_0_req_1); -- 
    cr_4384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(0), ack => type_cast_1418_inst_req_1); -- 
    cr_4320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(0), ack => type_cast_1402_inst_req_1); -- 
    rr_4226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(0), ack => ptr_deref_1382_load_0_req_0); -- 
    cr_4237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(0), ack => ptr_deref_1382_load_0_req_1); -- 
    cr_4256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(0), ack => type_cast_1386_inst_req_1); -- 
    rr_4290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(0), ack => ptr_deref_1398_load_0_req_0); -- 
    cr_4301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(0), ack => ptr_deref_1398_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_Sample/word_access_start/$exit
      -- CP-element group 1: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_Sample/word_access_start/word_0/ra
      -- 
    ra_4227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1382_load_0_ack_0, ack => sendOutput_CP_4163_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (12) 
      -- CP-element group 2: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_Update/word_access_complete/$exit
      -- CP-element group 2: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_Update/ptr_deref_1382_Merge/$entry
      -- CP-element group 2: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_Update/ptr_deref_1382_Merge/$exit
      -- CP-element group 2: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_Update/ptr_deref_1382_Merge/merge_req
      -- CP-element group 2: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1382_Update/ptr_deref_1382_Merge/merge_ack
      -- CP-element group 2: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1386_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1386_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1386_Sample/rr
      -- 
    ca_4238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1382_load_0_ack_1, ack => sendOutput_CP_4163_elements(2)); -- 
    rr_4251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(2), ack => type_cast_1386_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1386_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1386_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1386_Sample/ra
      -- 
    ra_4252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1386_inst_ack_0, ack => sendOutput_CP_4163_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	13 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1386_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1386_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1386_Update/ca
      -- 
    ca_4257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1386_inst_ack_1, ack => sendOutput_CP_4163_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_Sample/word_access_start/word_0/ra
      -- 
    ra_4291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1398_load_0_ack_0, ack => sendOutput_CP_4163_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (12) 
      -- CP-element group 6: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1402_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1402_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_Update/ptr_deref_1398_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_Update/ptr_deref_1398_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_Update/ptr_deref_1398_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1398_Update/ptr_deref_1398_Merge/merge_ack
      -- CP-element group 6: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1402_sample_start_
      -- 
    ca_4302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1398_load_0_ack_1, ack => sendOutput_CP_4163_elements(6)); -- 
    rr_4315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(6), ack => type_cast_1402_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1402_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1402_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1402_sample_completed_
      -- 
    ra_4316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1402_inst_ack_0, ack => sendOutput_CP_4163_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	13 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1402_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1402_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1402_update_completed_
      -- 
    ca_4321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1402_inst_ack_1, ack => sendOutput_CP_4163_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_Sample/word_access_start/word_0/ra
      -- 
    ra_4355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1414_load_0_ack_0, ack => sendOutput_CP_4163_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (12) 
      -- CP-element group 10: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_Update/ptr_deref_1414_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_Update/ptr_deref_1414_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1418_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1418_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_Update/ptr_deref_1414_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_Update/ptr_deref_1414_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1418_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/ptr_deref_1414_Update/word_access_complete/word_0/ca
      -- 
    ca_4366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1414_load_0_ack_1, ack => sendOutput_CP_4163_elements(10)); -- 
    rr_4379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(10), ack => type_cast_1418_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1418_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1418_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1418_Sample/$exit
      -- 
    ra_4380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1418_inst_ack_0, ack => sendOutput_CP_4163_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1418_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1418_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/type_cast_1418_Update/$exit
      -- 
    ca_4385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1418_inst_ack_1, ack => sendOutput_CP_4163_elements(12)); -- 
    -- CP-element group 13:  branch  join  transition  place  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: 	4 
    -- CP-element group 13: 	8 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (10) 
      -- CP-element group 13: 	 branch_block_stmt_1371/if_stmt_1436_if_link/$entry
      -- CP-element group 13: 	 branch_block_stmt_1371/if_stmt_1436_dead_link/$entry
      -- CP-element group 13: 	 branch_block_stmt_1371/if_stmt_1436_eval_test/$exit
      -- CP-element group 13: 	 branch_block_stmt_1371/if_stmt_1436_eval_test/branch_req
      -- CP-element group 13: 	 branch_block_stmt_1371/if_stmt_1436_else_link/$entry
      -- CP-element group 13: 	 branch_block_stmt_1371/R_cmp77_1437_place
      -- CP-element group 13: 	 branch_block_stmt_1371/if_stmt_1436_eval_test/$entry
      -- CP-element group 13: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435__exit__
      -- CP-element group 13: 	 branch_block_stmt_1371/if_stmt_1436__entry__
      -- CP-element group 13: 	 branch_block_stmt_1371/assign_stmt_1379_to_assign_stmt_1435/$exit
      -- 
    branch_req_4393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(13), ack => if_stmt_1436_branch_req_0); -- 
    sendOutput_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendOutput_CP_4163_elements(12) & sendOutput_CP_4163_elements(4) & sendOutput_CP_4163_elements(8);
      gj_sendOutput_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_4163_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (18) 
      -- CP-element group 14: 	 branch_block_stmt_1371/if_stmt_1436_if_link/if_choice_transition
      -- CP-element group 14: 	 branch_block_stmt_1371/merge_stmt_1442_PhiReqMerge
      -- CP-element group 14: 	 branch_block_stmt_1371/assign_stmt_1448_to_assign_stmt_1477/type_cast_1463_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1371/assign_stmt_1448_to_assign_stmt_1477/type_cast_1463_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1371/assign_stmt_1448_to_assign_stmt_1477/type_cast_1463_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1371/entry_bbx_xnph
      -- CP-element group 14: 	 branch_block_stmt_1371/assign_stmt_1448_to_assign_stmt_1477/type_cast_1463_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1371/assign_stmt_1448_to_assign_stmt_1477/type_cast_1463_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_1371/if_stmt_1436_if_link/$exit
      -- CP-element group 14: 	 branch_block_stmt_1371/assign_stmt_1448_to_assign_stmt_1477/type_cast_1463_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1371/assign_stmt_1448_to_assign_stmt_1477/$entry
      -- CP-element group 14: 	 branch_block_stmt_1371/merge_stmt_1442__exit__
      -- CP-element group 14: 	 branch_block_stmt_1371/assign_stmt_1448_to_assign_stmt_1477__entry__
      -- CP-element group 14: 	 branch_block_stmt_1371/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 14: 	 branch_block_stmt_1371/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 14: 	 branch_block_stmt_1371/merge_stmt_1442_PhiAck/$entry
      -- CP-element group 14: 	 branch_block_stmt_1371/merge_stmt_1442_PhiAck/$exit
      -- CP-element group 14: 	 branch_block_stmt_1371/merge_stmt_1442_PhiAck/dummy
      -- 
    if_choice_transition_4398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1436_branch_ack_1, ack => sendOutput_CP_4163_elements(14)); -- 
    rr_4415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(14), ack => type_cast_1463_inst_req_0); -- 
    cr_4420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(14), ack => type_cast_1463_inst_req_1); -- 
    -- CP-element group 15:  transition  place  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	72 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_1371/if_stmt_1436_else_link/$exit
      -- CP-element group 15: 	 branch_block_stmt_1371/entry_forx_xend
      -- CP-element group 15: 	 branch_block_stmt_1371/if_stmt_1436_else_link/else_choice_transition
      -- CP-element group 15: 	 branch_block_stmt_1371/entry_forx_xend_PhiReq/$entry
      -- CP-element group 15: 	 branch_block_stmt_1371/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_4402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1436_branch_ack_0, ack => sendOutput_CP_4163_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1371/assign_stmt_1448_to_assign_stmt_1477/type_cast_1463_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1371/assign_stmt_1448_to_assign_stmt_1477/type_cast_1463_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1371/assign_stmt_1448_to_assign_stmt_1477/type_cast_1463_Sample/ra
      -- 
    ra_4416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1463_inst_ack_0, ack => sendOutput_CP_4163_elements(16)); -- 
    -- CP-element group 17:  transition  place  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	66 
    -- CP-element group 17:  members (9) 
      -- CP-element group 17: 	 branch_block_stmt_1371/assign_stmt_1448_to_assign_stmt_1477/type_cast_1463_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1371/assign_stmt_1448_to_assign_stmt_1477/type_cast_1463_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1371/assign_stmt_1448_to_assign_stmt_1477/$exit
      -- CP-element group 17: 	 branch_block_stmt_1371/assign_stmt_1448_to_assign_stmt_1477/type_cast_1463_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1371/assign_stmt_1448_to_assign_stmt_1477__exit__
      -- CP-element group 17: 	 branch_block_stmt_1371/bbx_xnph_forx_xbody
      -- CP-element group 17: 	 branch_block_stmt_1371/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 17: 	 branch_block_stmt_1371/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1480/$entry
      -- CP-element group 17: 	 branch_block_stmt_1371/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1480/phi_stmt_1480_sources/$entry
      -- 
    ca_4421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1463_inst_ack_1, ack => sendOutput_CP_4163_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	71 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	63 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_final_index_sum_regn_Sample/ack
      -- CP-element group 18: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_final_index_sum_regn_sample_complete
      -- CP-element group 18: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_final_index_sum_regn_Sample/$exit
      -- 
    ack_4450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1492_index_offset_ack_0, ack => sendOutput_CP_4163_elements(18)); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	71 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (11) 
      -- CP-element group 19: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_root_address_calculated
      -- CP-element group 19: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_final_index_sum_regn_Update/ack
      -- CP-element group 19: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_base_plus_offset/$entry
      -- CP-element group 19: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_base_plus_offset/$exit
      -- CP-element group 19: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_base_plus_offset/sum_rename_req
      -- CP-element group 19: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_offset_calculated
      -- CP-element group 19: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/addr_of_1493_request/req
      -- CP-element group 19: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/addr_of_1493_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/addr_of_1493_request/$entry
      -- CP-element group 19: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_base_plus_offset/sum_rename_ack
      -- CP-element group 19: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_final_index_sum_regn_Update/$exit
      -- 
    ack_4455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1492_index_offset_ack_1, ack => sendOutput_CP_4163_elements(19)); -- 
    req_4464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(19), ack => addr_of_1493_final_reg_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/addr_of_1493_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/addr_of_1493_request/$exit
      -- CP-element group 20: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/addr_of_1493_request/ack
      -- 
    ack_4465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1493_final_reg_ack_0, ack => sendOutput_CP_4163_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	71 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (24) 
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/addr_of_1493_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_Sample/word_access_start/$entry
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_word_addrgen/$exit
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_base_addr_resize/base_resize_req
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_base_plus_offset/sum_rename_ack
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_word_addrgen/root_register_req
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_word_addrgen/$entry
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_base_addr_resize/$exit
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_root_address_calculated
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_base_plus_offset/$entry
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_word_address_calculated
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_Sample/word_access_start/word_0/rr
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_base_address_resized
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_base_addr_resize/base_resize_ack
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_base_plus_offset/sum_rename_req
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_base_address_calculated
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_base_plus_offset/$exit
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_base_addr_resize/$entry
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_Sample/word_access_start/word_0/$entry
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/addr_of_1493_complete/$exit
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_word_addrgen/root_register_ack
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/addr_of_1493_complete/ack
      -- CP-element group 21: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_Sample/$entry
      -- 
    ack_4470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1493_final_reg_ack_1, ack => sendOutput_CP_4163_elements(21)); -- 
    rr_4503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(21), ack => ptr_deref_1497_load_0_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (5) 
      -- CP-element group 22: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_Sample/word_access_start/word_0/ra
      -- CP-element group 22: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_Sample/word_access_start/$exit
      -- CP-element group 22: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_Sample/word_access_start/word_0/$exit
      -- 
    ra_4504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1497_load_0_ack_0, ack => sendOutput_CP_4163_elements(22)); -- 
    -- CP-element group 23:  fork  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	71 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	26 
    -- CP-element group 23: 	28 
    -- CP-element group 23: 	30 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	32 
    -- CP-element group 23: 	36 
    -- CP-element group 23: 	34 
    -- CP-element group 23: 	38 
    -- CP-element group 23:  members (33) 
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1531_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1511_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_Update/word_access_complete/$exit
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1521_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_Update/ptr_deref_1497_Merge/$entry
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1531_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1541_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1511_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1561_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1571_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_Update/ptr_deref_1497_Merge/merge_req
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1561_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1551_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1501_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1561_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1501_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1501_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1551_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1551_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_Update/word_access_complete/word_0/$exit
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1571_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1521_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1541_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1571_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_Update/ptr_deref_1497_Merge/merge_ack
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1541_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1511_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_Update/word_access_complete/word_0/ca
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1521_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_Update/ptr_deref_1497_Merge/$exit
      -- CP-element group 23: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1531_sample_start_
      -- 
    ca_4515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1497_load_0_ack_1, ack => sendOutput_CP_4163_elements(23)); -- 
    rr_4556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(23), ack => type_cast_1521_inst_req_0); -- 
    rr_4570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(23), ack => type_cast_1531_inst_req_0); -- 
    rr_4528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(23), ack => type_cast_1501_inst_req_0); -- 
    rr_4542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(23), ack => type_cast_1511_inst_req_0); -- 
    rr_4584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(23), ack => type_cast_1541_inst_req_0); -- 
    rr_4612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(23), ack => type_cast_1561_inst_req_0); -- 
    rr_4626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(23), ack => type_cast_1571_inst_req_0); -- 
    rr_4598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(23), ack => type_cast_1551_inst_req_0); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1501_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1501_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1501_sample_completed_
      -- 
    ra_4529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1501_inst_ack_0, ack => sendOutput_CP_4163_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	71 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	60 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1501_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1501_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1501_update_completed_
      -- 
    ca_4534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1501_inst_ack_1, ack => sendOutput_CP_4163_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	23 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1511_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1511_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1511_Sample/ra
      -- 
    ra_4543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1511_inst_ack_0, ack => sendOutput_CP_4163_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	71 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	57 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1511_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1511_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1511_Update/$exit
      -- 
    ca_4548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1511_inst_ack_1, ack => sendOutput_CP_4163_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	23 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1521_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1521_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1521_Sample/ra
      -- 
    ra_4557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1521_inst_ack_0, ack => sendOutput_CP_4163_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	71 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	54 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1521_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1521_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1521_Update/ca
      -- 
    ca_4562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1521_inst_ack_1, ack => sendOutput_CP_4163_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	23 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1531_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1531_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1531_Sample/ra
      -- 
    ra_4571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1531_inst_ack_0, ack => sendOutput_CP_4163_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	71 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	51 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1531_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1531_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1531_Update/$exit
      -- 
    ca_4576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1531_inst_ack_1, ack => sendOutput_CP_4163_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	23 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1541_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1541_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1541_sample_completed_
      -- 
    ra_4585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1541_inst_ack_0, ack => sendOutput_CP_4163_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	71 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	48 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1541_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1541_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1541_update_completed_
      -- 
    ca_4590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1541_inst_ack_1, ack => sendOutput_CP_4163_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1551_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1551_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1551_sample_completed_
      -- 
    ra_4599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1551_inst_ack_0, ack => sendOutput_CP_4163_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	71 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	45 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1551_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1551_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1551_Update/$exit
      -- 
    ca_4604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1551_inst_ack_1, ack => sendOutput_CP_4163_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	23 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1561_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1561_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1561_Sample/ra
      -- 
    ra_4613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1561_inst_ack_0, ack => sendOutput_CP_4163_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	71 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	42 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1561_Update/ca
      -- CP-element group 37: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1561_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1561_update_completed_
      -- 
    ca_4618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1561_inst_ack_1, ack => sendOutput_CP_4163_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	23 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1571_Sample/ra
      -- CP-element group 38: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1571_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1571_sample_completed_
      -- 
    ra_4627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1571_inst_ack_0, ack => sendOutput_CP_4163_elements(38)); -- 
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	71 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (6) 
      -- CP-element group 39: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1571_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1571_Update/ca
      -- CP-element group 39: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1571_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1573_Sample/req
      -- CP-element group 39: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1573_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1573_sample_start_
      -- 
    ca_4632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1571_inst_ack_1, ack => sendOutput_CP_4163_elements(39)); -- 
    req_4640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(39), ack => WPIPE_ConvTranspose_output_pipe_1573_inst_req_0); -- 
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (6) 
      -- CP-element group 40: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1573_Update/req
      -- CP-element group 40: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1573_Update/$entry
      -- CP-element group 40: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1573_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1573_update_start_
      -- CP-element group 40: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1573_Sample/ack
      -- CP-element group 40: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1573_Sample/$exit
      -- 
    ack_4641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1573_inst_ack_0, ack => sendOutput_CP_4163_elements(40)); -- 
    req_4645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(40), ack => WPIPE_ConvTranspose_output_pipe_1573_inst_req_1); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1573_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1573_Update/ack
      -- CP-element group 41: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1573_update_completed_
      -- 
    ack_4646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1573_inst_ack_1, ack => sendOutput_CP_4163_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	37 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1576_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1576_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1576_Sample/req
      -- 
    req_4654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(42), ack => WPIPE_ConvTranspose_output_pipe_1576_inst_req_0); -- 
    sendOutput_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_4163_elements(37) & sendOutput_CP_4163_elements(41);
      gj_sendOutput_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_4163_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1576_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1576_update_start_
      -- CP-element group 43: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1576_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1576_Sample/ack
      -- CP-element group 43: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1576_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1576_Update/req
      -- 
    ack_4655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1576_inst_ack_0, ack => sendOutput_CP_4163_elements(43)); -- 
    req_4659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(43), ack => WPIPE_ConvTranspose_output_pipe_1576_inst_req_1); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1576_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1576_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1576_Update/ack
      -- 
    ack_4660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1576_inst_ack_1, ack => sendOutput_CP_4163_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	35 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1579_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1579_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1579_Sample/req
      -- 
    req_4668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(45), ack => WPIPE_ConvTranspose_output_pipe_1579_inst_req_0); -- 
    sendOutput_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_4163_elements(35) & sendOutput_CP_4163_elements(44);
      gj_sendOutput_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_4163_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1579_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1579_update_start_
      -- CP-element group 46: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1579_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1579_Sample/ack
      -- CP-element group 46: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1579_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1579_Update/req
      -- 
    ack_4669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1579_inst_ack_0, ack => sendOutput_CP_4163_elements(46)); -- 
    req_4673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(46), ack => WPIPE_ConvTranspose_output_pipe_1579_inst_req_1); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1579_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1579_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1579_Update/ack
      -- 
    ack_4674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1579_inst_ack_1, ack => sendOutput_CP_4163_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	33 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1582_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1582_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1582_Sample/req
      -- 
    req_4682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(48), ack => WPIPE_ConvTranspose_output_pipe_1582_inst_req_0); -- 
    sendOutput_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_4163_elements(33) & sendOutput_CP_4163_elements(47);
      gj_sendOutput_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_4163_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1582_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1582_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1582_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1582_Sample/ack
      -- CP-element group 49: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1582_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1582_Update/req
      -- 
    ack_4683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1582_inst_ack_0, ack => sendOutput_CP_4163_elements(49)); -- 
    req_4687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(49), ack => WPIPE_ConvTranspose_output_pipe_1582_inst_req_1); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1582_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1582_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1582_Update/ack
      -- 
    ack_4688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1582_inst_ack_1, ack => sendOutput_CP_4163_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	31 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1585_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1585_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1585_Sample/req
      -- 
    req_4696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(51), ack => WPIPE_ConvTranspose_output_pipe_1585_inst_req_0); -- 
    sendOutput_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_4163_elements(31) & sendOutput_CP_4163_elements(50);
      gj_sendOutput_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_4163_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (6) 
      -- CP-element group 52: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1585_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1585_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1585_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1585_Sample/ack
      -- CP-element group 52: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1585_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1585_Update/req
      -- 
    ack_4697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1585_inst_ack_0, ack => sendOutput_CP_4163_elements(52)); -- 
    req_4701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(52), ack => WPIPE_ConvTranspose_output_pipe_1585_inst_req_1); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1585_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1585_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1585_Update/ack
      -- 
    ack_4702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1585_inst_ack_1, ack => sendOutput_CP_4163_elements(53)); -- 
    -- CP-element group 54:  join  transition  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	29 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1588_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1588_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1588_Sample/req
      -- 
    req_4710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(54), ack => WPIPE_ConvTranspose_output_pipe_1588_inst_req_0); -- 
    sendOutput_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_4163_elements(29) & sendOutput_CP_4163_elements(53);
      gj_sendOutput_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_4163_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (6) 
      -- CP-element group 55: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1588_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1588_update_start_
      -- CP-element group 55: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1588_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1588_Sample/ack
      -- CP-element group 55: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1588_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1588_Update/req
      -- 
    ack_4711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1588_inst_ack_0, ack => sendOutput_CP_4163_elements(55)); -- 
    req_4715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(55), ack => WPIPE_ConvTranspose_output_pipe_1588_inst_req_1); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1588_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1588_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1588_Update/ack
      -- 
    ack_4716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1588_inst_ack_1, ack => sendOutput_CP_4163_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	27 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1591_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1591_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1591_Sample/req
      -- 
    req_4724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(57), ack => WPIPE_ConvTranspose_output_pipe_1591_inst_req_0); -- 
    sendOutput_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_4163_elements(27) & sendOutput_CP_4163_elements(56);
      gj_sendOutput_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_4163_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (6) 
      -- CP-element group 58: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1591_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1591_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1591_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1591_Sample/ack
      -- CP-element group 58: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1591_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1591_Update/req
      -- 
    ack_4725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1591_inst_ack_0, ack => sendOutput_CP_4163_elements(58)); -- 
    req_4729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(58), ack => WPIPE_ConvTranspose_output_pipe_1591_inst_req_1); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1591_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1591_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1591_Update/ack
      -- 
    ack_4730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1591_inst_ack_1, ack => sendOutput_CP_4163_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	25 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1594_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1594_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1594_Sample/req
      -- 
    req_4738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(60), ack => WPIPE_ConvTranspose_output_pipe_1594_inst_req_0); -- 
    sendOutput_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_4163_elements(25) & sendOutput_CP_4163_elements(59);
      gj_sendOutput_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_4163_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1594_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1594_update_start_
      -- CP-element group 61: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1594_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1594_Sample/ack
      -- CP-element group 61: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1594_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1594_Update/req
      -- 
    ack_4739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1594_inst_ack_0, ack => sendOutput_CP_4163_elements(61)); -- 
    req_4743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(61), ack => WPIPE_ConvTranspose_output_pipe_1594_inst_req_1); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1594_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1594_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/WPIPE_ConvTranspose_output_pipe_1594_Update/ack
      -- 
    ack_4744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1594_inst_ack_1, ack => sendOutput_CP_4163_elements(62)); -- 
    -- CP-element group 63:  branch  join  transition  place  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	18 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (10) 
      -- CP-element group 63: 	 branch_block_stmt_1371/R_exitcond1_1609_place
      -- CP-element group 63: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/$exit
      -- CP-element group 63: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607__exit__
      -- CP-element group 63: 	 branch_block_stmt_1371/if_stmt_1608__entry__
      -- CP-element group 63: 	 branch_block_stmt_1371/if_stmt_1608_dead_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1371/if_stmt_1608_eval_test/$entry
      -- CP-element group 63: 	 branch_block_stmt_1371/if_stmt_1608_eval_test/$exit
      -- CP-element group 63: 	 branch_block_stmt_1371/if_stmt_1608_eval_test/branch_req
      -- CP-element group 63: 	 branch_block_stmt_1371/if_stmt_1608_if_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1371/if_stmt_1608_else_link/$entry
      -- 
    branch_req_4752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(63), ack => if_stmt_1608_branch_req_0); -- 
    sendOutput_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_4163_elements(18) & sendOutput_CP_4163_elements(62);
      gj_sendOutput_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_4163_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  merge  transition  place  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	72 
    -- CP-element group 64:  members (13) 
      -- CP-element group 64: 	 branch_block_stmt_1371/merge_stmt_1614_PhiReqMerge
      -- CP-element group 64: 	 branch_block_stmt_1371/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 64: 	 branch_block_stmt_1371/merge_stmt_1614__exit__
      -- CP-element group 64: 	 branch_block_stmt_1371/forx_xendx_xloopexit_forx_xend
      -- CP-element group 64: 	 branch_block_stmt_1371/if_stmt_1608_if_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_1371/if_stmt_1608_if_link/if_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_1371/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_1371/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 64: 	 branch_block_stmt_1371/merge_stmt_1614_PhiAck/$entry
      -- CP-element group 64: 	 branch_block_stmt_1371/merge_stmt_1614_PhiAck/$exit
      -- CP-element group 64: 	 branch_block_stmt_1371/merge_stmt_1614_PhiAck/dummy
      -- CP-element group 64: 	 branch_block_stmt_1371/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_1371/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_4757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1608_branch_ack_1, ack => sendOutput_CP_4163_elements(64)); -- 
    -- CP-element group 65:  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (12) 
      -- CP-element group 65: 	 branch_block_stmt_1371/forx_xbody_forx_xbody
      -- CP-element group 65: 	 branch_block_stmt_1371/if_stmt_1608_else_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_1371/if_stmt_1608_else_link/else_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_1371/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_1371/forx_xbody_forx_xbody_PhiReq/phi_stmt_1480/$entry
      -- CP-element group 65: 	 branch_block_stmt_1371/forx_xbody_forx_xbody_PhiReq/phi_stmt_1480/phi_stmt_1480_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_1371/forx_xbody_forx_xbody_PhiReq/phi_stmt_1480/phi_stmt_1480_sources/type_cast_1486/$entry
      -- CP-element group 65: 	 branch_block_stmt_1371/forx_xbody_forx_xbody_PhiReq/phi_stmt_1480/phi_stmt_1480_sources/type_cast_1486/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_1371/forx_xbody_forx_xbody_PhiReq/phi_stmt_1480/phi_stmt_1480_sources/type_cast_1486/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1371/forx_xbody_forx_xbody_PhiReq/phi_stmt_1480/phi_stmt_1480_sources/type_cast_1486/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_1371/forx_xbody_forx_xbody_PhiReq/phi_stmt_1480/phi_stmt_1480_sources/type_cast_1486/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1371/forx_xbody_forx_xbody_PhiReq/phi_stmt_1480/phi_stmt_1480_sources/type_cast_1486/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1608_branch_ack_0, ack => sendOutput_CP_4163_elements(65)); -- 
    rr_4805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(65), ack => type_cast_1486_inst_req_0); -- 
    cr_4810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(65), ack => type_cast_1486_inst_req_1); -- 
    -- CP-element group 66:  transition  output  delay-element  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	17 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	70 
    -- CP-element group 66:  members (5) 
      -- CP-element group 66: 	 branch_block_stmt_1371/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 66: 	 branch_block_stmt_1371/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1480/$exit
      -- CP-element group 66: 	 branch_block_stmt_1371/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1480/phi_stmt_1480_sources/$exit
      -- CP-element group 66: 	 branch_block_stmt_1371/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1480/phi_stmt_1480_sources/type_cast_1484_konst_delay_trans
      -- CP-element group 66: 	 branch_block_stmt_1371/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1480/phi_stmt_1480_req
      -- 
    phi_stmt_1480_req_4786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1480_req_4786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(66), ack => phi_stmt_1480_req_0); -- 
    -- Element group sendOutput_CP_4163_elements(66) is a control-delay.
    cp_element_66_delay: control_delay_element  generic map(name => " 66_delay", delay_value => 1)  port map(req => sendOutput_CP_4163_elements(17), ack => sendOutput_CP_4163_elements(66), clk => clk, reset =>reset);
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_1371/forx_xbody_forx_xbody_PhiReq/phi_stmt_1480/phi_stmt_1480_sources/type_cast_1486/SplitProtocol/Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_1371/forx_xbody_forx_xbody_PhiReq/phi_stmt_1480/phi_stmt_1480_sources/type_cast_1486/SplitProtocol/Sample/ra
      -- 
    ra_4806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1486_inst_ack_0, ack => sendOutput_CP_4163_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	65 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1371/forx_xbody_forx_xbody_PhiReq/phi_stmt_1480/phi_stmt_1480_sources/type_cast_1486/SplitProtocol/Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_1371/forx_xbody_forx_xbody_PhiReq/phi_stmt_1480/phi_stmt_1480_sources/type_cast_1486/SplitProtocol/Update/ca
      -- 
    ca_4811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1486_inst_ack_1, ack => sendOutput_CP_4163_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (6) 
      -- CP-element group 69: 	 branch_block_stmt_1371/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1371/forx_xbody_forx_xbody_PhiReq/phi_stmt_1480/$exit
      -- CP-element group 69: 	 branch_block_stmt_1371/forx_xbody_forx_xbody_PhiReq/phi_stmt_1480/phi_stmt_1480_sources/$exit
      -- CP-element group 69: 	 branch_block_stmt_1371/forx_xbody_forx_xbody_PhiReq/phi_stmt_1480/phi_stmt_1480_sources/type_cast_1486/$exit
      -- CP-element group 69: 	 branch_block_stmt_1371/forx_xbody_forx_xbody_PhiReq/phi_stmt_1480/phi_stmt_1480_sources/type_cast_1486/SplitProtocol/$exit
      -- CP-element group 69: 	 branch_block_stmt_1371/forx_xbody_forx_xbody_PhiReq/phi_stmt_1480/phi_stmt_1480_req
      -- 
    phi_stmt_1480_req_4812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1480_req_4812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(69), ack => phi_stmt_1480_req_1); -- 
    sendOutput_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_4163_elements(67) & sendOutput_CP_4163_elements(68);
      gj_sendOutput_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_4163_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  merge  transition  place  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	66 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_1371/merge_stmt_1479_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_1371/merge_stmt_1479_PhiAck/$entry
      -- 
    sendOutput_CP_4163_elements(70) <= OrReduce(sendOutput_CP_4163_elements(66) & sendOutput_CP_4163_elements(69));
    -- CP-element group 71:  fork  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	27 
    -- CP-element group 71: 	29 
    -- CP-element group 71: 	18 
    -- CP-element group 71: 	19 
    -- CP-element group 71: 	21 
    -- CP-element group 71: 	23 
    -- CP-element group 71: 	25 
    -- CP-element group 71: 	31 
    -- CP-element group 71: 	37 
    -- CP-element group 71: 	33 
    -- CP-element group 71: 	35 
    -- CP-element group 71: 	39 
    -- CP-element group 71:  members (53) 
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_index_resized_1
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_final_index_sum_regn_Update/req
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_Update/word_access_complete/$entry
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_index_scale_1/$entry
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1531_update_start_
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1531_Update/cr
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/addr_of_1493_update_start_
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_index_scale_1/$exit
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_update_start_
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1521_Update/cr
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_index_resize_1/index_resize_req
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_final_index_sum_regn_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1511_Update/cr
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1521_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_final_index_sum_regn_Sample/req
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1501_Update/cr
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_Update/word_access_complete/word_0/$entry
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1501_update_start_
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1501_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_index_resize_1/$exit
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_index_scale_1/scale_rename_ack
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1571_Update/cr
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_index_resize_1/$entry
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1551_update_start_
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/$entry
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1571_update_start_
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_final_index_sum_regn_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1571_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1551_Update/cr
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1511_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1561_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1511_update_start_
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1561_update_start_
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_index_resize_1/index_resize_ack
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1521_update_start_
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1541_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_final_index_sum_regn_update_start
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1541_Update/cr
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1561_Update/cr
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_index_computed_1
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1541_update_start_
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/ptr_deref_1497_Update/word_access_complete/word_0/cr
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1551_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/addr_of_1493_complete/$entry
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_index_scale_1/scale_rename_req
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/array_obj_ref_1492_index_scaled_1
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/type_cast_1531_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607/addr_of_1493_complete/req
      -- CP-element group 71: 	 branch_block_stmt_1371/merge_stmt_1479__exit__
      -- CP-element group 71: 	 branch_block_stmt_1371/assign_stmt_1494_to_assign_stmt_1607__entry__
      -- CP-element group 71: 	 branch_block_stmt_1371/merge_stmt_1479_PhiAck/$exit
      -- CP-element group 71: 	 branch_block_stmt_1371/merge_stmt_1479_PhiAck/phi_stmt_1480_ack
      -- 
    phi_stmt_1480_ack_4817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1480_ack_0, ack => sendOutput_CP_4163_elements(71)); -- 
    req_4454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(71), ack => array_obj_ref_1492_index_offset_req_1); -- 
    cr_4575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(71), ack => type_cast_1531_inst_req_1); -- 
    cr_4561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(71), ack => type_cast_1521_inst_req_1); -- 
    cr_4547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(71), ack => type_cast_1511_inst_req_1); -- 
    req_4449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(71), ack => array_obj_ref_1492_index_offset_req_0); -- 
    cr_4533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(71), ack => type_cast_1501_inst_req_1); -- 
    cr_4631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(71), ack => type_cast_1571_inst_req_1); -- 
    cr_4603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(71), ack => type_cast_1551_inst_req_1); -- 
    cr_4589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(71), ack => type_cast_1541_inst_req_1); -- 
    cr_4617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(71), ack => type_cast_1561_inst_req_1); -- 
    cr_4514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(71), ack => ptr_deref_1497_load_0_req_1); -- 
    req_4469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_4163_elements(71), ack => addr_of_1493_final_reg_req_1); -- 
    -- CP-element group 72:  merge  transition  place  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	15 
    -- CP-element group 72: 	64 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (16) 
      -- CP-element group 72: 	 $exit
      -- CP-element group 72: 	 branch_block_stmt_1371/$exit
      -- CP-element group 72: 	 branch_block_stmt_1371/branch_block_stmt_1371__exit__
      -- CP-element group 72: 	 branch_block_stmt_1371/merge_stmt_1616__exit__
      -- CP-element group 72: 	 branch_block_stmt_1371/return__
      -- CP-element group 72: 	 branch_block_stmt_1371/merge_stmt_1618__exit__
      -- CP-element group 72: 	 branch_block_stmt_1371/merge_stmt_1616_PhiReqMerge
      -- CP-element group 72: 	 branch_block_stmt_1371/merge_stmt_1616_PhiAck/$entry
      -- CP-element group 72: 	 branch_block_stmt_1371/merge_stmt_1616_PhiAck/$exit
      -- CP-element group 72: 	 branch_block_stmt_1371/merge_stmt_1616_PhiAck/dummy
      -- CP-element group 72: 	 branch_block_stmt_1371/return___PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_1371/return___PhiReq/$exit
      -- CP-element group 72: 	 branch_block_stmt_1371/merge_stmt_1618_PhiReqMerge
      -- CP-element group 72: 	 branch_block_stmt_1371/merge_stmt_1618_PhiAck/$entry
      -- CP-element group 72: 	 branch_block_stmt_1371/merge_stmt_1618_PhiAck/$exit
      -- CP-element group 72: 	 branch_block_stmt_1371/merge_stmt_1618_PhiAck/dummy
      -- 
    sendOutput_CP_4163_elements(72) <= OrReduce(sendOutput_CP_4163_elements(15) & sendOutput_CP_4163_elements(64));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar_1491_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1491_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_1492_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1492_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1492_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1492_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1492_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1492_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_1494 : std_logic_vector(31 downto 0);
    signal cmp77_1435 : std_logic_vector(0 downto 0);
    signal conv15_1502 : std_logic_vector(7 downto 0);
    signal conv21_1512 : std_logic_vector(7 downto 0);
    signal conv27_1522 : std_logic_vector(7 downto 0);
    signal conv2_1403 : std_logic_vector(31 downto 0);
    signal conv33_1532 : std_logic_vector(7 downto 0);
    signal conv39_1542 : std_logic_vector(7 downto 0);
    signal conv45_1552 : std_logic_vector(7 downto 0);
    signal conv4_1419 : std_logic_vector(31 downto 0);
    signal conv51_1562 : std_logic_vector(7 downto 0);
    signal conv57_1572 : std_logic_vector(7 downto 0);
    signal conv_1387 : std_logic_vector(31 downto 0);
    signal exitcond1_1607 : std_logic_vector(0 downto 0);
    signal iNsTr_0_1379 : std_logic_vector(31 downto 0);
    signal iNsTr_1_1395 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1411 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1464 : std_logic_vector(63 downto 0);
    signal indvar_1480 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1602 : std_logic_vector(63 downto 0);
    signal mul5_1429 : std_logic_vector(31 downto 0);
    signal mul_1424 : std_logic_vector(31 downto 0);
    signal ptr_deref_1382_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1382_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1382_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1382_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1382_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1398_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1398_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1398_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1398_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1398_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1414_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1414_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1414_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1414_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1414_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1497_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1497_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1497_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1497_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1497_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr18_1508 : std_logic_vector(63 downto 0);
    signal shr24_1518 : std_logic_vector(63 downto 0);
    signal shr30_1528 : std_logic_vector(63 downto 0);
    signal shr36_1538 : std_logic_vector(63 downto 0);
    signal shr42_1548 : std_logic_vector(63 downto 0);
    signal shr48_1558 : std_logic_vector(63 downto 0);
    signal shr54_1568 : std_logic_vector(63 downto 0);
    signal tmp12_1498 : std_logic_vector(63 downto 0);
    signal tmp1_1399 : std_logic_vector(15 downto 0);
    signal tmp3_1415 : std_logic_vector(15 downto 0);
    signal tmp84_1448 : std_logic_vector(31 downto 0);
    signal tmp84x_xop_1460 : std_logic_vector(31 downto 0);
    signal tmp85_1454 : std_logic_vector(0 downto 0);
    signal tmp88_1477 : std_logic_vector(63 downto 0);
    signal tmp_1383 : std_logic_vector(15 downto 0);
    signal type_cast_1433_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1446_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1452_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1458_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1468_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1475_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1484_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1486_wire : std_logic_vector(63 downto 0);
    signal type_cast_1506_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1516_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1526_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1536_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1546_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1556_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1566_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1600_wire_constant : std_logic_vector(63 downto 0);
    signal xx_xop_1470 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1492_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1492_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1492_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1492_resized_base_address <= "00000000000000";
    iNsTr_0_1379 <= "00000000000000000000000000000100";
    iNsTr_1_1395 <= "00000000000000000000000000000101";
    iNsTr_2_1411 <= "00000000000000000000000000000110";
    ptr_deref_1382_word_offset_0 <= "0000000";
    ptr_deref_1398_word_offset_0 <= "0000000";
    ptr_deref_1414_word_offset_0 <= "0000000";
    ptr_deref_1497_word_offset_0 <= "00000000000000";
    type_cast_1433_wire_constant <= "00000000000000000000000000000011";
    type_cast_1446_wire_constant <= "00000000000000000000000000000010";
    type_cast_1452_wire_constant <= "00000000000000000000000000000001";
    type_cast_1458_wire_constant <= "11111111111111111111111111111111";
    type_cast_1468_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1475_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1484_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1506_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1516_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1526_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1536_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1546_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1556_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1566_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1600_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_1480: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1484_wire_constant & type_cast_1486_wire;
      req <= phi_stmt_1480_req_0 & phi_stmt_1480_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1480",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1480_ack_0,
          idata => idata,
          odata => indvar_1480,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1480
    -- flow-through select operator MUX_1476_inst
    tmp88_1477 <= xx_xop_1470 when (tmp85_1454(0) /=  '0') else type_cast_1475_wire_constant;
    addr_of_1493_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1493_final_reg_req_0;
      addr_of_1493_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1493_final_reg_req_1;
      addr_of_1493_final_reg_ack_1<= rack(0);
      addr_of_1493_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1493_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1492_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1494,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1386_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1386_inst_req_0;
      type_cast_1386_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1386_inst_req_1;
      type_cast_1386_inst_ack_1<= rack(0);
      type_cast_1386_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1386_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_1383,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1387,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1402_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1402_inst_req_0;
      type_cast_1402_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1402_inst_req_1;
      type_cast_1402_inst_ack_1<= rack(0);
      type_cast_1402_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1402_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1_1399,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2_1403,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1418_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1418_inst_req_0;
      type_cast_1418_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1418_inst_req_1;
      type_cast_1418_inst_ack_1<= rack(0);
      type_cast_1418_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1418_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3_1415,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_1419,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1463_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1463_inst_req_0;
      type_cast_1463_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1463_inst_req_1;
      type_cast_1463_inst_ack_1<= rack(0);
      type_cast_1463_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1463_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp84x_xop_1460,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_4_1464,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1486_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1486_inst_req_0;
      type_cast_1486_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1486_inst_req_1;
      type_cast_1486_inst_ack_1<= rack(0);
      type_cast_1486_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1486_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1602,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1486_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1501_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1501_inst_req_0;
      type_cast_1501_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1501_inst_req_1;
      type_cast_1501_inst_ack_1<= rack(0);
      type_cast_1501_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1501_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp12_1498,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv15_1502,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1511_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1511_inst_req_0;
      type_cast_1511_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1511_inst_req_1;
      type_cast_1511_inst_ack_1<= rack(0);
      type_cast_1511_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1511_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr18_1508,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv21_1512,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1521_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1521_inst_req_0;
      type_cast_1521_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1521_inst_req_1;
      type_cast_1521_inst_ack_1<= rack(0);
      type_cast_1521_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1521_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr24_1518,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv27_1522,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1531_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1531_inst_req_0;
      type_cast_1531_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1531_inst_req_1;
      type_cast_1531_inst_ack_1<= rack(0);
      type_cast_1531_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1531_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr30_1528,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv33_1532,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1541_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1541_inst_req_0;
      type_cast_1541_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1541_inst_req_1;
      type_cast_1541_inst_ack_1<= rack(0);
      type_cast_1541_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1541_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr36_1538,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_1542,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1551_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1551_inst_req_0;
      type_cast_1551_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1551_inst_req_1;
      type_cast_1551_inst_ack_1<= rack(0);
      type_cast_1551_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1551_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr42_1548,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv45_1552,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1561_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1561_inst_req_0;
      type_cast_1561_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1561_inst_req_1;
      type_cast_1561_inst_ack_1<= rack(0);
      type_cast_1561_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1561_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr48_1558,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv51_1562,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1571_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1571_inst_req_0;
      type_cast_1571_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1571_inst_req_1;
      type_cast_1571_inst_ack_1<= rack(0);
      type_cast_1571_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1571_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr54_1568,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv57_1572,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1492_index_1_rename
    process(R_indvar_1491_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1491_resized;
      ov(13 downto 0) := iv;
      R_indvar_1491_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1492_index_1_resize
    process(indvar_1480) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1480;
      ov := iv(13 downto 0);
      R_indvar_1491_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1492_root_address_inst
    process(array_obj_ref_1492_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1492_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1492_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1382_addr_0
    process(ptr_deref_1382_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1382_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1382_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1382_base_resize
    process(iNsTr_0_1379) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_1379;
      ov := iv(6 downto 0);
      ptr_deref_1382_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1382_gather_scatter
    process(ptr_deref_1382_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1382_data_0;
      ov(15 downto 0) := iv;
      tmp_1383 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1382_root_address_inst
    process(ptr_deref_1382_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1382_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1382_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1398_addr_0
    process(ptr_deref_1398_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1398_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1398_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1398_base_resize
    process(iNsTr_1_1395) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_1_1395;
      ov := iv(6 downto 0);
      ptr_deref_1398_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1398_gather_scatter
    process(ptr_deref_1398_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1398_data_0;
      ov(15 downto 0) := iv;
      tmp1_1399 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1398_root_address_inst
    process(ptr_deref_1398_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1398_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1398_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1414_addr_0
    process(ptr_deref_1414_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1414_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1414_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1414_base_resize
    process(iNsTr_2_1411) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1411;
      ov := iv(6 downto 0);
      ptr_deref_1414_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1414_gather_scatter
    process(ptr_deref_1414_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1414_data_0;
      ov(15 downto 0) := iv;
      tmp3_1415 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1414_root_address_inst
    process(ptr_deref_1414_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1414_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1414_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1497_addr_0
    process(ptr_deref_1497_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1497_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1497_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1497_base_resize
    process(arrayidx_1494) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1494;
      ov := iv(13 downto 0);
      ptr_deref_1497_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1497_gather_scatter
    process(ptr_deref_1497_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1497_data_0;
      ov(63 downto 0) := iv;
      tmp12_1498 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1497_root_address_inst
    process(ptr_deref_1497_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1497_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1497_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1436_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp77_1435;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1436_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1436_branch_req_0,
          ack0 => if_stmt_1436_branch_ack_0,
          ack1 => if_stmt_1436_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1608_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1607;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1608_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1608_branch_req_0,
          ack0 => if_stmt_1608_branch_ack_0,
          ack1 => if_stmt_1608_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1459_inst
    process(tmp84_1448) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp84_1448, type_cast_1458_wire_constant, tmp_var);
      tmp84x_xop_1460 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1469_inst
    process(iNsTr_4_1464) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_4_1464, type_cast_1468_wire_constant, tmp_var);
      xx_xop_1470 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1601_inst
    process(indvar_1480) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1480, type_cast_1600_wire_constant, tmp_var);
      indvarx_xnext_1602 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1606_inst
    process(indvarx_xnext_1602, tmp88_1477) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1602, tmp88_1477, tmp_var);
      exitcond1_1607 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1447_inst
    process(mul5_1429) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul5_1429, type_cast_1446_wire_constant, tmp_var);
      tmp84_1448 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1507_inst
    process(tmp12_1498) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp12_1498, type_cast_1506_wire_constant, tmp_var);
      shr18_1508 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1517_inst
    process(tmp12_1498) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp12_1498, type_cast_1516_wire_constant, tmp_var);
      shr24_1518 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1527_inst
    process(tmp12_1498) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp12_1498, type_cast_1526_wire_constant, tmp_var);
      shr30_1528 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1537_inst
    process(tmp12_1498) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp12_1498, type_cast_1536_wire_constant, tmp_var);
      shr36_1538 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1547_inst
    process(tmp12_1498) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp12_1498, type_cast_1546_wire_constant, tmp_var);
      shr42_1548 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1557_inst
    process(tmp12_1498) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp12_1498, type_cast_1556_wire_constant, tmp_var);
      shr48_1558 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1567_inst
    process(tmp12_1498) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp12_1498, type_cast_1566_wire_constant, tmp_var);
      shr54_1568 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1423_inst
    process(conv2_1403, conv_1387) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv2_1403, conv_1387, tmp_var);
      mul_1424 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1428_inst
    process(mul_1424, conv4_1419) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_1424, conv4_1419, tmp_var);
      mul5_1429 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1434_inst
    process(mul5_1429) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul5_1429, type_cast_1433_wire_constant, tmp_var);
      cmp77_1435 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1453_inst
    process(tmp84_1448) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp84_1448, type_cast_1452_wire_constant, tmp_var);
      tmp85_1454 <= tmp_var; --
    end process;
    -- shared split operator group (16) : array_obj_ref_1492_index_offset 
    ApIntAdd_group_16: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1491_scaled;
      array_obj_ref_1492_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1492_index_offset_req_0;
      array_obj_ref_1492_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1492_index_offset_req_1;
      array_obj_ref_1492_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_16_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_16_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared load operator group (0) : ptr_deref_1382_load_0 ptr_deref_1398_load_0 ptr_deref_1414_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1382_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1398_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1414_load_0_req_0;
      ptr_deref_1382_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1398_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1414_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1382_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1398_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1414_load_0_req_1;
      ptr_deref_1382_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1398_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1414_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1382_word_address_0 & ptr_deref_1398_word_address_0 & ptr_deref_1414_word_address_0;
      ptr_deref_1382_data_0 <= data_out(47 downto 32);
      ptr_deref_1398_data_0 <= data_out(31 downto 16);
      ptr_deref_1414_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(15 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1497_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1497_load_0_req_0;
      ptr_deref_1497_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1497_load_0_req_1;
      ptr_deref_1497_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1497_word_address_0;
      ptr_deref_1497_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(13 downto 0),
          mtag => memory_space_6_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(63 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared outport operator group (0) : WPIPE_ConvTranspose_output_pipe_1573_inst WPIPE_ConvTranspose_output_pipe_1576_inst WPIPE_ConvTranspose_output_pipe_1579_inst WPIPE_ConvTranspose_output_pipe_1582_inst WPIPE_ConvTranspose_output_pipe_1585_inst WPIPE_ConvTranspose_output_pipe_1588_inst WPIPE_ConvTranspose_output_pipe_1591_inst WPIPE_ConvTranspose_output_pipe_1594_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1573_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1576_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1579_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1582_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1585_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1588_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1591_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1594_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1573_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1576_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1579_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1582_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1585_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1588_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1591_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1594_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1573_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1576_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1579_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1582_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1585_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1588_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1591_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1594_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1573_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1576_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1579_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1582_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1585_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1588_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1591_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1594_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv57_1572 & conv51_1562 & conv45_1552 & conv39_1542 & conv33_1532 & conv27_1522 & conv21_1512 & conv15_1502;
      ConvTranspose_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendOutput_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity testConfigure is -- 
  generic (tag_length : integer); 
  port ( -- 
    ret_val_x_x : out  std_logic_vector(15 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_7_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_8_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity testConfigure;
architecture testConfigure_arch of testConfigure is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 16)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ret_val_x_x_buffer :  std_logic_vector(15 downto 0);
  signal testConfigure_CP_0_start: Boolean;
  signal testConfigure_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_711_load_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_364_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_364_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_506_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_845_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_506_inst_ack_0 : boolean;
  signal ptr_deref_711_load_0_req_0 : boolean;
  signal ptr_deref_496_store_0_ack_1 : boolean;
  signal array_obj_ref_841_index_offset_req_0 : boolean;
  signal ptr_deref_496_store_0_ack_0 : boolean;
  signal ptr_deref_496_store_0_req_0 : boolean;
  signal ptr_deref_496_store_0_req_1 : boolean;
  signal type_cast_916_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_894_inst_req_1 : boolean;
  signal if_stmt_770_branch_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_36_inst_ack_1 : boolean;
  signal ptr_deref_392_store_0_ack_1 : boolean;
  signal addr_of_389_final_reg_ack_1 : boolean;
  signal ptr_deref_392_store_0_req_1 : boolean;
  signal type_cast_368_inst_ack_1 : boolean;
  signal ptr_deref_392_store_0_ack_0 : boolean;
  signal type_cast_368_inst_req_1 : boolean;
  signal ptr_deref_392_store_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_36_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_36_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_36_inst_req_1 : boolean;
  signal array_obj_ref_841_index_offset_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_912_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_481_inst_req_1 : boolean;
  signal type_cast_40_inst_req_0 : boolean;
  signal type_cast_40_inst_ack_0 : boolean;
  signal type_cast_40_inst_req_1 : boolean;
  signal type_cast_40_inst_ack_1 : boolean;
  signal if_stmt_436_branch_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_418_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_418_inst_req_0 : boolean;
  signal ptr_deref_49_store_0_req_0 : boolean;
  signal ptr_deref_49_store_0_ack_0 : boolean;
  signal ptr_deref_49_store_0_req_1 : boolean;
  signal ptr_deref_49_store_0_ack_1 : boolean;
  signal type_cast_457_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_ack_0 : boolean;
  signal addr_of_389_final_reg_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_ack_1 : boolean;
  signal type_cast_63_inst_req_0 : boolean;
  signal type_cast_63_inst_ack_0 : boolean;
  signal type_cast_63_inst_req_1 : boolean;
  signal type_cast_63_inst_ack_1 : boolean;
  signal array_obj_ref_841_index_offset_ack_1 : boolean;
  signal ptr_deref_77_store_0_req_0 : boolean;
  signal ptr_deref_77_store_0_ack_0 : boolean;
  signal type_cast_368_inst_ack_0 : boolean;
  signal ptr_deref_77_store_0_req_1 : boolean;
  signal ptr_deref_77_store_0_ack_1 : boolean;
  signal if_stmt_785_branch_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_88_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_88_inst_ack_0 : boolean;
  signal addr_of_389_final_reg_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_88_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_88_inst_ack_1 : boolean;
  signal type_cast_1222_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_481_inst_ack_1 : boolean;
  signal if_stmt_785_branch_ack_1 : boolean;
  signal type_cast_92_inst_req_0 : boolean;
  signal type_cast_92_inst_ack_0 : boolean;
  signal type_cast_92_inst_req_1 : boolean;
  signal type_cast_92_inst_ack_1 : boolean;
  signal type_cast_368_inst_req_0 : boolean;
  signal if_stmt_94_branch_req_0 : boolean;
  signal type_cast_457_inst_req_1 : boolean;
  signal if_stmt_94_branch_ack_1 : boolean;
  signal if_stmt_94_branch_ack_0 : boolean;
  signal type_cast_125_inst_req_0 : boolean;
  signal type_cast_125_inst_ack_0 : boolean;
  signal type_cast_125_inst_req_1 : boolean;
  signal type_cast_125_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_466_inst_ack_1 : boolean;
  signal type_cast_285_inst_ack_0 : boolean;
  signal type_cast_285_inst_req_1 : boolean;
  signal type_cast_285_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_402_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_402_inst_req_0 : boolean;
  signal array_obj_ref_131_index_offset_req_0 : boolean;
  signal array_obj_ref_131_index_offset_ack_0 : boolean;
  signal addr_of_389_final_reg_req_0 : boolean;
  signal array_obj_ref_131_index_offset_req_1 : boolean;
  signal array_obj_ref_131_index_offset_ack_1 : boolean;
  signal type_cast_485_inst_ack_0 : boolean;
  signal if_stmt_785_branch_ack_0 : boolean;
  signal addr_of_132_final_reg_req_0 : boolean;
  signal addr_of_132_final_reg_ack_0 : boolean;
  signal addr_of_132_final_reg_req_1 : boolean;
  signal addr_of_132_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_466_inst_req_1 : boolean;
  signal type_cast_406_inst_ack_1 : boolean;
  signal ptr_deref_135_store_0_req_0 : boolean;
  signal ptr_deref_135_store_0_ack_0 : boolean;
  signal ptr_deref_135_store_0_req_1 : boolean;
  signal type_cast_406_inst_req_1 : boolean;
  signal ptr_deref_135_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_145_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_145_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_145_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_145_inst_ack_1 : boolean;
  signal STORE_padding_477_store_0_ack_1 : boolean;
  signal STORE_padding_477_store_0_req_1 : boolean;
  signal type_cast_422_inst_ack_1 : boolean;
  signal STORE_padding_452_store_0_ack_1 : boolean;
  signal type_cast_149_inst_req_0 : boolean;
  signal type_cast_149_inst_ack_0 : boolean;
  signal type_cast_149_inst_req_1 : boolean;
  signal type_cast_149_inst_ack_1 : boolean;
  signal if_stmt_770_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_466_inst_ack_0 : boolean;
  signal type_cast_422_inst_req_1 : boolean;
  signal type_cast_862_inst_req_0 : boolean;
  signal ptr_deref_414_store_0_ack_1 : boolean;
  signal type_cast_406_inst_ack_0 : boolean;
  signal STORE_padding_452_store_0_req_1 : boolean;
  signal ptr_deref_414_store_0_req_1 : boolean;
  signal ptr_deref_157_store_0_req_0 : boolean;
  signal ptr_deref_157_store_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_845_inst_ack_1 : boolean;
  signal ptr_deref_157_store_0_req_1 : boolean;
  signal type_cast_406_inst_req_0 : boolean;
  signal ptr_deref_157_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_466_inst_req_0 : boolean;
  signal type_cast_422_inst_ack_0 : boolean;
  signal type_cast_422_inst_req_0 : boolean;
  signal ptr_deref_1332_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_894_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_481_inst_ack_0 : boolean;
  signal type_cast_470_inst_ack_1 : boolean;
  signal ptr_deref_174_load_0_req_0 : boolean;
  signal ptr_deref_174_load_0_ack_0 : boolean;
  signal ptr_deref_174_load_0_req_1 : boolean;
  signal ptr_deref_174_load_0_ack_1 : boolean;
  signal type_cast_880_inst_ack_0 : boolean;
  signal type_cast_178_inst_req_0 : boolean;
  signal type_cast_178_inst_ack_0 : boolean;
  signal type_cast_178_inst_req_1 : boolean;
  signal type_cast_178_inst_ack_1 : boolean;
  signal type_cast_485_inst_req_0 : boolean;
  signal type_cast_470_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_189_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_189_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_189_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_189_inst_ack_1 : boolean;
  signal array_obj_ref_841_index_offset_ack_0 : boolean;
  signal type_cast_862_inst_ack_0 : boolean;
  signal type_cast_193_inst_req_0 : boolean;
  signal type_cast_193_inst_ack_0 : boolean;
  signal type_cast_193_inst_req_1 : boolean;
  signal type_cast_193_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_481_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_364_inst_ack_1 : boolean;
  signal if_stmt_195_branch_req_0 : boolean;
  signal type_cast_457_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_364_inst_req_1 : boolean;
  signal if_stmt_195_branch_ack_1 : boolean;
  signal if_stmt_195_branch_ack_0 : boolean;
  signal if_stmt_436_branch_ack_0 : boolean;
  signal ptr_deref_414_store_0_ack_0 : boolean;
  signal ptr_deref_414_store_0_req_0 : boolean;
  signal type_cast_470_inst_ack_0 : boolean;
  signal ptr_deref_223_store_0_req_0 : boolean;
  signal ptr_deref_223_store_0_ack_0 : boolean;
  signal type_cast_470_inst_req_0 : boolean;
  signal ptr_deref_223_store_0_req_1 : boolean;
  signal ptr_deref_223_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_233_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_233_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_233_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_233_inst_ack_1 : boolean;
  signal type_cast_485_inst_ack_1 : boolean;
  signal type_cast_457_inst_req_0 : boolean;
  signal STORE_padding_477_store_0_ack_0 : boolean;
  signal type_cast_812_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_876_inst_req_1 : boolean;
  signal STORE_padding_452_store_0_ack_0 : boolean;
  signal type_cast_237_inst_req_0 : boolean;
  signal type_cast_237_inst_ack_0 : boolean;
  signal type_cast_731_inst_ack_1 : boolean;
  signal type_cast_237_inst_req_1 : boolean;
  signal type_cast_237_inst_ack_1 : boolean;
  signal if_stmt_354_branch_ack_0 : boolean;
  signal STORE_padding_452_store_0_req_0 : boolean;
  signal ptr_deref_251_store_0_req_0 : boolean;
  signal ptr_deref_251_store_0_ack_0 : boolean;
  signal ptr_deref_251_store_0_req_1 : boolean;
  signal ptr_deref_251_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_402_inst_ack_1 : boolean;
  signal if_stmt_436_branch_ack_1 : boolean;
  signal if_stmt_260_branch_req_0 : boolean;
  signal type_cast_812_inst_ack_0 : boolean;
  signal ptr_deref_711_load_0_req_1 : boolean;
  signal if_stmt_260_branch_ack_1 : boolean;
  signal if_stmt_354_branch_ack_1 : boolean;
  signal if_stmt_260_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_402_inst_req_1 : boolean;
  signal type_cast_285_inst_req_0 : boolean;
  signal array_obj_ref_291_index_offset_req_0 : boolean;
  signal array_obj_ref_291_index_offset_ack_0 : boolean;
  signal array_obj_ref_291_index_offset_req_1 : boolean;
  signal array_obj_ref_291_index_offset_ack_1 : boolean;
  signal STORE_padding_477_store_0_req_0 : boolean;
  signal ptr_deref_1332_store_0_req_1 : boolean;
  signal addr_of_292_final_reg_req_0 : boolean;
  signal addr_of_292_final_reg_ack_0 : boolean;
  signal addr_of_292_final_reg_req_1 : boolean;
  signal addr_of_292_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_418_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_418_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_295_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_295_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_295_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_295_inst_ack_1 : boolean;
  signal type_cast_485_inst_req_1 : boolean;
  signal type_cast_299_inst_req_0 : boolean;
  signal type_cast_299_inst_ack_0 : boolean;
  signal type_cast_299_inst_req_1 : boolean;
  signal type_cast_299_inst_ack_1 : boolean;
  signal type_cast_812_inst_req_1 : boolean;
  signal type_cast_812_inst_ack_1 : boolean;
  signal type_cast_731_inst_req_0 : boolean;
  signal ptr_deref_302_store_0_req_0 : boolean;
  signal ptr_deref_302_store_0_ack_0 : boolean;
  signal ptr_deref_711_load_0_ack_1 : boolean;
  signal type_cast_731_inst_ack_0 : boolean;
  signal ptr_deref_302_store_0_req_1 : boolean;
  signal ptr_deref_302_store_0_ack_1 : boolean;
  signal type_cast_862_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_312_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_312_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_312_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_312_inst_ack_1 : boolean;
  signal type_cast_316_inst_req_0 : boolean;
  signal type_cast_316_inst_ack_0 : boolean;
  signal type_cast_880_inst_req_0 : boolean;
  signal type_cast_316_inst_req_1 : boolean;
  signal type_cast_316_inst_ack_1 : boolean;
  signal type_cast_731_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_876_inst_ack_1 : boolean;
  signal ptr_deref_324_store_0_req_0 : boolean;
  signal ptr_deref_324_store_0_ack_0 : boolean;
  signal ptr_deref_324_store_0_req_1 : boolean;
  signal ptr_deref_324_store_0_ack_1 : boolean;
  signal ptr_deref_341_load_0_req_0 : boolean;
  signal ptr_deref_341_load_0_ack_0 : boolean;
  signal ptr_deref_341_load_0_req_1 : boolean;
  signal ptr_deref_341_load_0_ack_1 : boolean;
  signal type_cast_345_inst_req_0 : boolean;
  signal type_cast_345_inst_ack_0 : boolean;
  signal type_cast_345_inst_req_1 : boolean;
  signal type_cast_345_inst_ack_1 : boolean;
  signal if_stmt_354_branch_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_506_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_506_inst_ack_1 : boolean;
  signal type_cast_113_inst_ack_1 : boolean;
  signal type_cast_880_inst_ack_1 : boolean;
  signal if_stmt_770_branch_req_0 : boolean;
  signal type_cast_510_inst_req_0 : boolean;
  signal type_cast_510_inst_ack_0 : boolean;
  signal type_cast_510_inst_req_1 : boolean;
  signal type_cast_510_inst_ack_1 : boolean;
  signal type_cast_916_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_845_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_845_inst_req_0 : boolean;
  signal ptr_deref_526_store_0_req_0 : boolean;
  signal ptr_deref_526_store_0_ack_0 : boolean;
  signal ptr_deref_526_store_0_req_1 : boolean;
  signal ptr_deref_526_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_894_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_530_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_530_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_530_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_530_inst_ack_1 : boolean;
  signal type_cast_898_inst_ack_1 : boolean;
  signal type_cast_205_inst_req_1 : boolean;
  signal type_cast_898_inst_req_1 : boolean;
  signal type_cast_1222_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_858_inst_ack_1 : boolean;
  signal type_cast_534_inst_req_0 : boolean;
  signal type_cast_1222_inst_req_1 : boolean;
  signal type_cast_534_inst_ack_0 : boolean;
  signal type_cast_534_inst_req_1 : boolean;
  signal type_cast_534_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_894_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_858_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_858_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_912_inst_ack_0 : boolean;
  signal ptr_deref_727_load_0_ack_1 : boolean;
  signal ptr_deref_545_store_0_req_0 : boolean;
  signal type_cast_747_inst_ack_1 : boolean;
  signal ptr_deref_545_store_0_ack_0 : boolean;
  signal ptr_deref_727_load_0_req_1 : boolean;
  signal ptr_deref_545_store_0_req_1 : boolean;
  signal type_cast_747_inst_req_1 : boolean;
  signal ptr_deref_545_store_0_ack_1 : boolean;
  signal type_cast_916_inst_ack_0 : boolean;
  signal type_cast_113_inst_req_1 : boolean;
  signal type_cast_699_inst_ack_1 : boolean;
  signal type_cast_115_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_555_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_555_inst_ack_0 : boolean;
  signal type_cast_715_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_555_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_555_inst_ack_1 : boolean;
  signal type_cast_898_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_912_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_858_inst_req_0 : boolean;
  signal type_cast_747_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_876_inst_ack_0 : boolean;
  signal type_cast_559_inst_req_0 : boolean;
  signal if_stmt_1199_branch_req_0 : boolean;
  signal type_cast_559_inst_ack_0 : boolean;
  signal type_cast_559_inst_req_1 : boolean;
  signal type_cast_559_inst_ack_1 : boolean;
  signal type_cast_916_inst_req_0 : boolean;
  signal type_cast_747_inst_req_0 : boolean;
  signal array_obj_ref_1328_index_offset_req_0 : boolean;
  signal ptr_deref_575_store_0_req_0 : boolean;
  signal ptr_deref_575_store_0_ack_0 : boolean;
  signal ptr_deref_575_store_0_req_1 : boolean;
  signal ptr_deref_575_store_0_ack_1 : boolean;
  signal type_cast_898_inst_req_0 : boolean;
  signal type_cast_205_inst_req_0 : boolean;
  signal type_cast_715_inst_req_1 : boolean;
  signal type_cast_115_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_579_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_579_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_579_inst_req_1 : boolean;
  signal array_obj_ref_1328_index_offset_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_579_inst_ack_1 : boolean;
  signal type_cast_880_inst_req_1 : boolean;
  signal type_cast_583_inst_req_0 : boolean;
  signal type_cast_583_inst_ack_0 : boolean;
  signal type_cast_583_inst_req_1 : boolean;
  signal type_cast_583_inst_ack_1 : boolean;
  signal addr_of_842_final_reg_ack_1 : boolean;
  signal if_stmt_1347_branch_req_0 : boolean;
  signal addr_of_842_final_reg_req_1 : boolean;
  signal ptr_deref_743_load_0_ack_1 : boolean;
  signal type_cast_1222_inst_ack_1 : boolean;
  signal ptr_deref_594_store_0_req_0 : boolean;
  signal ptr_deref_743_load_0_req_1 : boolean;
  signal ptr_deref_594_store_0_ack_0 : boolean;
  signal ptr_deref_594_store_0_req_1 : boolean;
  signal ptr_deref_594_store_0_ack_1 : boolean;
  signal type_cast_699_inst_req_1 : boolean;
  signal type_cast_862_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_604_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_604_inst_ack_0 : boolean;
  signal type_cast_715_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_604_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_604_inst_ack_1 : boolean;
  signal if_stmt_1347_branch_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_876_inst_req_0 : boolean;
  signal type_cast_608_inst_req_0 : boolean;
  signal type_cast_608_inst_ack_0 : boolean;
  signal phi_stmt_110_req_0 : boolean;
  signal type_cast_608_inst_req_1 : boolean;
  signal addr_of_842_final_reg_ack_0 : boolean;
  signal type_cast_608_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_912_inst_ack_1 : boolean;
  signal type_cast_849_inst_ack_1 : boolean;
  signal type_cast_849_inst_req_1 : boolean;
  signal type_cast_849_inst_ack_0 : boolean;
  signal addr_of_842_final_reg_req_0 : boolean;
  signal type_cast_715_inst_req_0 : boolean;
  signal ptr_deref_743_load_0_ack_0 : boolean;
  signal ptr_deref_743_load_0_req_0 : boolean;
  signal array_obj_ref_1328_index_offset_req_1 : boolean;
  signal ptr_deref_727_load_0_ack_0 : boolean;
  signal ptr_deref_727_load_0_req_0 : boolean;
  signal ptr_deref_624_store_0_req_0 : boolean;
  signal ptr_deref_624_store_0_ack_0 : boolean;
  signal ptr_deref_624_store_0_req_1 : boolean;
  signal ptr_deref_624_store_0_ack_1 : boolean;
  signal type_cast_699_inst_ack_0 : boolean;
  signal array_obj_ref_1328_index_offset_ack_1 : boolean;
  signal type_cast_699_inst_req_0 : boolean;
  signal ptr_deref_637_load_0_req_0 : boolean;
  signal ptr_deref_637_load_0_ack_0 : boolean;
  signal ptr_deref_637_load_0_req_1 : boolean;
  signal ptr_deref_637_load_0_ack_1 : boolean;
  signal type_cast_849_inst_req_0 : boolean;
  signal type_cast_641_inst_req_0 : boolean;
  signal type_cast_641_inst_ack_0 : boolean;
  signal type_cast_641_inst_req_1 : boolean;
  signal type_cast_641_inst_ack_1 : boolean;
  signal ptr_deref_653_load_0_req_0 : boolean;
  signal ptr_deref_653_load_0_ack_0 : boolean;
  signal ptr_deref_653_load_0_req_1 : boolean;
  signal ptr_deref_653_load_0_ack_1 : boolean;
  signal if_stmt_1347_branch_ack_0 : boolean;
  signal type_cast_657_inst_req_0 : boolean;
  signal type_cast_657_inst_ack_0 : boolean;
  signal type_cast_657_inst_req_1 : boolean;
  signal type_cast_657_inst_ack_1 : boolean;
  signal if_stmt_1199_branch_ack_1 : boolean;
  signal ptr_deref_1250_load_0_req_1 : boolean;
  signal ptr_deref_669_load_0_req_0 : boolean;
  signal ptr_deref_669_load_0_ack_0 : boolean;
  signal ptr_deref_669_load_0_req_1 : boolean;
  signal ptr_deref_669_load_0_ack_1 : boolean;
  signal type_cast_673_inst_req_0 : boolean;
  signal type_cast_673_inst_ack_0 : boolean;
  signal type_cast_673_inst_req_1 : boolean;
  signal type_cast_673_inst_ack_1 : boolean;
  signal ptr_deref_695_load_0_req_0 : boolean;
  signal ptr_deref_695_load_0_ack_0 : boolean;
  signal ptr_deref_695_load_0_req_1 : boolean;
  signal ptr_deref_695_load_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_930_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_930_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_930_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_930_inst_ack_1 : boolean;
  signal type_cast_212_inst_req_1 : boolean;
  signal type_cast_205_inst_ack_0 : boolean;
  signal type_cast_1238_inst_ack_1 : boolean;
  signal type_cast_934_inst_req_0 : boolean;
  signal type_cast_934_inst_ack_0 : boolean;
  signal type_cast_934_inst_req_1 : boolean;
  signal type_cast_934_inst_ack_1 : boolean;
  signal ptr_deref_1332_store_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_948_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_948_inst_ack_0 : boolean;
  signal ptr_deref_1218_load_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_948_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_948_inst_ack_1 : boolean;
  signal ptr_deref_1332_store_0_req_0 : boolean;
  signal type_cast_1238_inst_req_1 : boolean;
  signal phi_stmt_110_ack_0 : boolean;
  signal type_cast_952_inst_req_0 : boolean;
  signal type_cast_952_inst_ack_0 : boolean;
  signal type_cast_113_inst_ack_0 : boolean;
  signal type_cast_952_inst_req_1 : boolean;
  signal type_cast_952_inst_ack_1 : boolean;
  signal ptr_deref_1218_load_0_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_966_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_966_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_966_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_966_inst_ack_1 : boolean;
  signal type_cast_1238_inst_ack_0 : boolean;
  signal type_cast_115_inst_ack_1 : boolean;
  signal type_cast_970_inst_req_0 : boolean;
  signal type_cast_970_inst_ack_0 : boolean;
  signal type_cast_113_inst_req_0 : boolean;
  signal type_cast_970_inst_req_1 : boolean;
  signal type_cast_970_inst_ack_1 : boolean;
  signal type_cast_1238_inst_req_0 : boolean;
  signal type_cast_1299_inst_ack_1 : boolean;
  signal type_cast_1299_inst_req_1 : boolean;
  signal ptr_deref_978_store_0_req_0 : boolean;
  signal ptr_deref_978_store_0_ack_0 : boolean;
  signal ptr_deref_978_store_0_req_1 : boolean;
  signal ptr_deref_978_store_0_ack_1 : boolean;
  signal if_stmt_992_branch_req_0 : boolean;
  signal if_stmt_992_branch_ack_1 : boolean;
  signal ptr_deref_1250_load_0_ack_0 : boolean;
  signal if_stmt_992_branch_ack_0 : boolean;
  signal ptr_deref_1250_load_0_req_0 : boolean;
  signal if_stmt_1199_branch_ack_0 : boolean;
  signal type_cast_115_inst_req_1 : boolean;
  signal type_cast_1019_inst_req_0 : boolean;
  signal type_cast_1019_inst_ack_0 : boolean;
  signal type_cast_1019_inst_req_1 : boolean;
  signal type_cast_1299_inst_ack_0 : boolean;
  signal type_cast_1019_inst_ack_1 : boolean;
  signal phi_stmt_103_req_0 : boolean;
  signal phi_stmt_103_ack_0 : boolean;
  signal type_cast_106_inst_ack_1 : boolean;
  signal type_cast_106_inst_req_1 : boolean;
  signal array_obj_ref_1048_index_offset_req_0 : boolean;
  signal type_cast_1299_inst_req_0 : boolean;
  signal array_obj_ref_1048_index_offset_ack_0 : boolean;
  signal array_obj_ref_1048_index_offset_req_1 : boolean;
  signal array_obj_ref_1048_index_offset_ack_1 : boolean;
  signal ptr_deref_1234_load_0_ack_1 : boolean;
  signal addr_of_1049_final_reg_req_0 : boolean;
  signal addr_of_1049_final_reg_ack_0 : boolean;
  signal addr_of_1049_final_reg_req_1 : boolean;
  signal addr_of_1049_final_reg_ack_1 : boolean;
  signal phi_stmt_209_req_0 : boolean;
  signal type_cast_106_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1052_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1052_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1052_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1052_inst_ack_1 : boolean;
  signal ptr_deref_1234_load_0_req_1 : boolean;
  signal type_cast_1056_inst_req_0 : boolean;
  signal type_cast_1056_inst_ack_0 : boolean;
  signal type_cast_1056_inst_req_1 : boolean;
  signal if_stmt_1272_branch_ack_0 : boolean;
  signal type_cast_1056_inst_ack_1 : boolean;
  signal type_cast_106_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1065_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1065_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1065_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1065_inst_ack_1 : boolean;
  signal type_cast_212_inst_ack_0 : boolean;
  signal phi_stmt_202_req_0 : boolean;
  signal type_cast_1069_inst_req_0 : boolean;
  signal if_stmt_1272_branch_ack_1 : boolean;
  signal type_cast_1069_inst_ack_0 : boolean;
  signal type_cast_1069_inst_req_1 : boolean;
  signal type_cast_1069_inst_ack_1 : boolean;
  signal type_cast_212_inst_ack_1 : boolean;
  signal ptr_deref_1218_load_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1083_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1083_inst_ack_0 : boolean;
  signal ptr_deref_1218_load_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1083_inst_req_1 : boolean;
  signal if_stmt_1272_branch_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1083_inst_ack_1 : boolean;
  signal type_cast_212_inst_req_0 : boolean;
  signal type_cast_1087_inst_req_0 : boolean;
  signal type_cast_1087_inst_ack_0 : boolean;
  signal type_cast_1087_inst_req_1 : boolean;
  signal type_cast_1087_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1101_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1101_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1101_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1101_inst_ack_1 : boolean;
  signal type_cast_205_inst_ack_1 : boolean;
  signal ptr_deref_1234_load_0_ack_0 : boolean;
  signal phi_stmt_103_req_1 : boolean;
  signal type_cast_1105_inst_req_0 : boolean;
  signal type_cast_1105_inst_ack_0 : boolean;
  signal type_cast_1105_inst_req_1 : boolean;
  signal type_cast_1254_inst_ack_1 : boolean;
  signal type_cast_1105_inst_ack_1 : boolean;
  signal phi_stmt_202_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1119_inst_req_0 : boolean;
  signal type_cast_1254_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1119_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1119_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1119_inst_ack_1 : boolean;
  signal ptr_deref_1234_load_0_req_0 : boolean;
  signal phi_stmt_110_req_1 : boolean;
  signal type_cast_1123_inst_req_0 : boolean;
  signal type_cast_1123_inst_ack_0 : boolean;
  signal type_cast_1123_inst_req_1 : boolean;
  signal type_cast_1254_inst_ack_0 : boolean;
  signal type_cast_1123_inst_ack_1 : boolean;
  signal addr_of_1329_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1137_inst_req_0 : boolean;
  signal type_cast_1254_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1137_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1137_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1137_inst_ack_1 : boolean;
  signal type_cast_1141_inst_req_0 : boolean;
  signal type_cast_1141_inst_ack_0 : boolean;
  signal type_cast_1141_inst_req_1 : boolean;
  signal type_cast_1141_inst_ack_1 : boolean;
  signal addr_of_1329_final_reg_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1155_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1155_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1155_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1155_inst_ack_1 : boolean;
  signal type_cast_1159_inst_req_0 : boolean;
  signal type_cast_1159_inst_ack_0 : boolean;
  signal type_cast_1159_inst_req_1 : boolean;
  signal type_cast_1159_inst_ack_1 : boolean;
  signal addr_of_1329_final_reg_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1173_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1173_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1173_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_1173_inst_ack_1 : boolean;
  signal type_cast_1177_inst_req_0 : boolean;
  signal type_cast_1177_inst_ack_0 : boolean;
  signal type_cast_1177_inst_req_1 : boolean;
  signal ptr_deref_1250_load_0_ack_1 : boolean;
  signal type_cast_1177_inst_ack_1 : boolean;
  signal addr_of_1329_final_reg_req_0 : boolean;
  signal ptr_deref_1185_store_0_req_0 : boolean;
  signal ptr_deref_1185_store_0_ack_0 : boolean;
  signal ptr_deref_1185_store_0_req_1 : boolean;
  signal ptr_deref_1185_store_0_ack_1 : boolean;
  signal type_cast_214_inst_req_0 : boolean;
  signal type_cast_214_inst_ack_0 : boolean;
  signal type_cast_214_inst_req_1 : boolean;
  signal type_cast_214_inst_ack_1 : boolean;
  signal phi_stmt_209_req_1 : boolean;
  signal phi_stmt_209_ack_0 : boolean;
  signal type_cast_272_inst_req_0 : boolean;
  signal type_cast_272_inst_ack_0 : boolean;
  signal type_cast_272_inst_req_1 : boolean;
  signal type_cast_272_inst_ack_1 : boolean;
  signal phi_stmt_269_req_0 : boolean;
  signal phi_stmt_269_req_1 : boolean;
  signal phi_stmt_269_ack_0 : boolean;
  signal phi_stmt_372_req_0 : boolean;
  signal type_cast_382_inst_req_0 : boolean;
  signal type_cast_382_inst_ack_0 : boolean;
  signal type_cast_382_inst_req_1 : boolean;
  signal type_cast_382_inst_ack_1 : boolean;
  signal phi_stmt_379_req_0 : boolean;
  signal type_cast_378_inst_req_0 : boolean;
  signal type_cast_378_inst_ack_0 : boolean;
  signal type_cast_378_inst_req_1 : boolean;
  signal type_cast_378_inst_ack_1 : boolean;
  signal phi_stmt_372_req_1 : boolean;
  signal type_cast_384_inst_req_0 : boolean;
  signal type_cast_384_inst_ack_0 : boolean;
  signal type_cast_384_inst_req_1 : boolean;
  signal type_cast_384_inst_ack_1 : boolean;
  signal phi_stmt_379_req_1 : boolean;
  signal phi_stmt_372_ack_0 : boolean;
  signal phi_stmt_379_ack_0 : boolean;
  signal type_cast_446_inst_req_0 : boolean;
  signal type_cast_446_inst_ack_0 : boolean;
  signal type_cast_446_inst_req_1 : boolean;
  signal type_cast_446_inst_ack_1 : boolean;
  signal phi_stmt_443_req_0 : boolean;
  signal type_cast_450_inst_req_0 : boolean;
  signal type_cast_450_inst_ack_0 : boolean;
  signal type_cast_450_inst_req_1 : boolean;
  signal type_cast_450_inst_ack_1 : boolean;
  signal phi_stmt_447_req_0 : boolean;
  signal phi_stmt_443_ack_0 : boolean;
  signal phi_stmt_447_ack_0 : boolean;
  signal phi_stmt_829_req_0 : boolean;
  signal type_cast_835_inst_req_0 : boolean;
  signal type_cast_835_inst_ack_0 : boolean;
  signal type_cast_835_inst_req_1 : boolean;
  signal type_cast_835_inst_ack_1 : boolean;
  signal phi_stmt_829_req_1 : boolean;
  signal phi_stmt_829_ack_0 : boolean;
  signal phi_stmt_1036_req_0 : boolean;
  signal type_cast_1042_inst_req_0 : boolean;
  signal type_cast_1042_inst_ack_0 : boolean;
  signal type_cast_1042_inst_req_1 : boolean;
  signal type_cast_1042_inst_ack_1 : boolean;
  signal phi_stmt_1036_req_1 : boolean;
  signal phi_stmt_1036_ack_0 : boolean;
  signal phi_stmt_1316_req_0 : boolean;
  signal type_cast_1322_inst_req_0 : boolean;
  signal type_cast_1322_inst_ack_0 : boolean;
  signal type_cast_1322_inst_req_1 : boolean;
  signal type_cast_1322_inst_ack_1 : boolean;
  signal phi_stmt_1316_req_1 : boolean;
  signal phi_stmt_1316_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "testConfigure_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  testConfigure_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "testConfigure_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 16) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  ret_val_x_x_buffer <= "0000000000000001";
  out_buffer_data_in(15 downto 0) <= ret_val_x_x_buffer;
  ret_val_x_x <= out_buffer_data_out(15 downto 0);
  out_buffer_data_in(tag_length + 15 downto 16) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 15 downto 16);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= testConfigure_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  testConfigure_CP_0: Block -- control-path 
    signal testConfigure_CP_0_elements: BooleanArray(408 downto 0);
    -- 
  begin -- 
    testConfigure_CP_0_elements(0) <= testConfigure_CP_0_start;
    testConfigure_CP_0_symbol <= testConfigure_CP_0_elements(408);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	15 
    -- CP-element group 0: 	19 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (59) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_34/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/branch_block_stmt_34__entry__
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93__entry__
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_36_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_36_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_36_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_40_update_start_
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_40_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_40_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_update_start_
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_63_update_start_
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_63_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_63_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_update_start_
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_92_update_start_
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_92_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_92_Update/cr
      -- 
    rr_118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => RPIPE_ConvTranspose_input_pipe_36_inst_req_0); -- 
    cr_137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => type_cast_40_inst_req_1); -- 
    cr_187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => ptr_deref_49_store_0_req_1); -- 
    cr_215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => type_cast_63_inst_req_1); -- 
    cr_265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => ptr_deref_77_store_0_req_1); -- 
    cr_293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => type_cast_92_inst_req_1); -- 
    -- CP-element group 1:  merge  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	386 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	119 
    -- CP-element group 1:  members (2) 
      -- CP-element group 1: 	 branch_block_stmt_34/merge_stmt_442__exit__
      -- CP-element group 1: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769__entry__
      -- 
    testConfigure_CP_0_elements(1) <= testConfigure_CP_0_elements(386);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_36_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_36_update_start_
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_36_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_36_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_36_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_36_Update/cr
      -- 
    ra_119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_36_inst_ack_0, ack => testConfigure_CP_0_elements(2)); -- 
    cr_123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(2), ack => RPIPE_ConvTranspose_input_pipe_36_inst_req_1); -- 
    -- CP-element group 3:  fork  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	9 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_36_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_40_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_36_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_36_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_40_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_40_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_59_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_59_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_59_Sample/rr
      -- 
    ca_124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_36_inst_ack_1, ack => testConfigure_CP_0_elements(3)); -- 
    rr_196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(3), ack => RPIPE_ConvTranspose_input_pipe_59_inst_req_0); -- 
    rr_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(3), ack => type_cast_40_inst_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_40_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_40_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_40_Sample/ra
      -- 
    ra_133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_40_inst_ack_0, ack => testConfigure_CP_0_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_40_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_40_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_40_Update/ca
      -- 
    ca_138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_40_inst_ack_1, ack => testConfigure_CP_0_elements(5)); -- 
    -- CP-element group 6:  join  transition  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_Sample/ptr_deref_49_Split/$entry
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_Sample/ptr_deref_49_Split/$exit
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_Sample/ptr_deref_49_Split/split_req
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_Sample/ptr_deref_49_Split/split_ack
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_Sample/word_access_start/$entry
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_Sample/word_access_start/word_0/$entry
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_Sample/word_access_start/word_0/rr
      -- 
    rr_176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(6), ack => ptr_deref_49_store_0_req_0); -- 
    testConfigure_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "testConfigure_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(0) & testConfigure_CP_0_elements(5);
      gj_testConfigure_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	20 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_Sample/word_access_start/word_0/ra
      -- 
    ra_177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_49_store_0_ack_0, ack => testConfigure_CP_0_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_Update/word_access_complete/word_0/ca
      -- 
    ca_188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_49_store_0_ack_1, ack => testConfigure_CP_0_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	3 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_59_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_59_update_start_
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_59_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_59_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_59_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_59_Update/cr
      -- 
    ra_197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_59_inst_ack_0, ack => testConfigure_CP_0_elements(9)); -- 
    cr_201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(9), ack => RPIPE_ConvTranspose_input_pipe_59_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	16 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_59_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_59_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_59_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_63_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_63_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_63_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_88_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_88_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_88_Sample/rr
      -- 
    ca_202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_59_inst_ack_1, ack => testConfigure_CP_0_elements(10)); -- 
    rr_274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(10), ack => RPIPE_ConvTranspose_input_pipe_88_inst_req_0); -- 
    rr_210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(10), ack => type_cast_63_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_63_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_63_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_63_Sample/ra
      -- 
    ra_211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_63_inst_ack_0, ack => testConfigure_CP_0_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_63_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_63_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_63_Update/ca
      -- 
    ca_216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_63_inst_ack_1, ack => testConfigure_CP_0_elements(12)); -- 
    -- CP-element group 13:  join  transition  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: 	20 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (9) 
      -- CP-element group 13: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_Sample/ptr_deref_77_Split/$entry
      -- CP-element group 13: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_Sample/ptr_deref_77_Split/$exit
      -- CP-element group 13: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_Sample/ptr_deref_77_Split/split_req
      -- CP-element group 13: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_Sample/ptr_deref_77_Split/split_ack
      -- CP-element group 13: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_Sample/word_access_start/$entry
      -- CP-element group 13: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_Sample/word_access_start/word_0/$entry
      -- CP-element group 13: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_Sample/word_access_start/word_0/rr
      -- 
    rr_254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(13), ack => ptr_deref_77_store_0_req_0); -- 
    testConfigure_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(0) & testConfigure_CP_0_elements(20) & testConfigure_CP_0_elements(12);
      gj_testConfigure_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (5) 
      -- CP-element group 14: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_Sample/word_access_start/$exit
      -- CP-element group 14: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_Sample/word_access_start/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_Sample/word_access_start/word_0/ra
      -- 
    ra_255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_77_store_0_ack_0, ack => testConfigure_CP_0_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	0 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	21 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_Update/word_access_complete/$exit
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_Update/word_access_complete/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_77_Update/word_access_complete/word_0/ca
      -- 
    ca_266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_77_store_0_ack_1, ack => testConfigure_CP_0_elements(15)); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	10 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_88_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_88_update_start_
      -- CP-element group 16: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_88_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_88_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_88_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_88_Update/cr
      -- 
    ra_275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_88_inst_ack_0, ack => testConfigure_CP_0_elements(16)); -- 
    cr_279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(16), ack => RPIPE_ConvTranspose_input_pipe_88_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_88_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_88_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/RPIPE_ConvTranspose_input_pipe_88_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_92_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_92_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_92_Sample/rr
      -- 
    ca_280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_88_inst_ack_1, ack => testConfigure_CP_0_elements(17)); -- 
    rr_288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(17), ack => type_cast_92_inst_req_0); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_92_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_92_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_92_Sample/ra
      -- 
    ra_289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_92_inst_ack_0, ack => testConfigure_CP_0_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	0 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_92_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_92_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/type_cast_92_Update/ca
      -- 
    ca_294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_92_inst_ack_1, ack => testConfigure_CP_0_elements(19)); -- 
    -- CP-element group 20:  transition  delay-element  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	7 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	13 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/ptr_deref_49_ptr_deref_77_delay
      -- 
    -- Element group testConfigure_CP_0_elements(20) is a control-delay.
    cp_element_20_delay: control_delay_element  generic map(name => " 20_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(7), ack => testConfigure_CP_0_elements(20), clk => clk, reset =>reset);
    -- CP-element group 21:  branch  join  transition  place  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: 	15 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (10) 
      -- CP-element group 21: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93__exit__
      -- CP-element group 21: 	 branch_block_stmt_34/if_stmt_94__entry__
      -- CP-element group 21: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_93/$exit
      -- CP-element group 21: 	 branch_block_stmt_34/if_stmt_94_dead_link/$entry
      -- CP-element group 21: 	 branch_block_stmt_34/if_stmt_94_eval_test/$entry
      -- CP-element group 21: 	 branch_block_stmt_34/if_stmt_94_eval_test/$exit
      -- CP-element group 21: 	 branch_block_stmt_34/if_stmt_94_eval_test/branch_req
      -- CP-element group 21: 	 branch_block_stmt_34/R_cmp316_95_place
      -- CP-element group 21: 	 branch_block_stmt_34/if_stmt_94_if_link/$entry
      -- CP-element group 21: 	 branch_block_stmt_34/if_stmt_94_else_link/$entry
      -- 
    branch_req_303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(21), ack => if_stmt_94_branch_req_0); -- 
    testConfigure_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(8) & testConfigure_CP_0_elements(15) & testConfigure_CP_0_elements(19);
      gj_testConfigure_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  fork  transition  place  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	346 
    -- CP-element group 22: 	347 
    -- CP-element group 22:  members (12) 
      -- CP-element group 22: 	 branch_block_stmt_34/if_stmt_94_if_link/$exit
      -- CP-element group 22: 	 branch_block_stmt_34/if_stmt_94_if_link/if_choice_transition
      -- CP-element group 22: 	 branch_block_stmt_34/entry_forx_xend
      -- CP-element group 22: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_212/SplitProtocol/Update/cr
      -- CP-element group 22: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/$entry
      -- CP-element group 22: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_212/$entry
      -- CP-element group 22: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_209/$entry
      -- CP-element group 22: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_212/SplitProtocol/Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_212/SplitProtocol/Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_212/SplitProtocol/Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/$entry
      -- CP-element group 22: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_212/SplitProtocol/$entry
      -- 
    if_choice_transition_308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_94_branch_ack_1, ack => testConfigure_CP_0_elements(22)); -- 
    cr_3626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(22), ack => type_cast_212_inst_req_1); -- 
    rr_3621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(22), ack => type_cast_212_inst_req_0); -- 
    -- CP-element group 23:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	333 
    -- CP-element group 23: 	334 
    -- CP-element group 23: 	335 
    -- CP-element group 23:  members (22) 
      -- CP-element group 23: 	 branch_block_stmt_34/merge_stmt_100__exit__
      -- CP-element group 23: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody
      -- CP-element group 23: 	 branch_block_stmt_34/merge_stmt_100_PhiReqMerge
      -- CP-element group 23: 	 branch_block_stmt_34/if_stmt_94_else_link/$exit
      -- CP-element group 23: 	 branch_block_stmt_34/if_stmt_94_else_link/else_choice_transition
      -- CP-element group 23: 	 branch_block_stmt_34/entry_forx_xbodyx_xpreheader
      -- CP-element group 23: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_113/SplitProtocol/Update/cr
      -- CP-element group 23: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_113/SplitProtocol/Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_113/SplitProtocol/Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_113/SplitProtocol/Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_113/SplitProtocol/$entry
      -- CP-element group 23: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_103/$entry
      -- CP-element group 23: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/$entry
      -- CP-element group 23: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_113/$entry
      -- CP-element group 23: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/$entry
      -- CP-element group 23: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_110/$entry
      -- CP-element group 23: 	 branch_block_stmt_34/merge_stmt_100_PhiAck/dummy
      -- CP-element group 23: 	 branch_block_stmt_34/merge_stmt_100_PhiAck/$exit
      -- CP-element group 23: 	 branch_block_stmt_34/merge_stmt_100_PhiAck/$entry
      -- CP-element group 23: 	 branch_block_stmt_34/entry_forx_xbodyx_xpreheader_PhiReq/$exit
      -- CP-element group 23: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_103/phi_stmt_103_sources/$entry
      -- CP-element group 23: 	 branch_block_stmt_34/entry_forx_xbodyx_xpreheader_PhiReq/$entry
      -- 
    else_choice_transition_312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_94_branch_ack_0, ack => testConfigure_CP_0_elements(23)); -- 
    cr_3559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(23), ack => type_cast_113_inst_req_1); -- 
    rr_3554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(23), ack => type_cast_113_inst_req_0); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	341 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_125_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_125_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_125_Sample/ra
      -- 
    ra_326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_125_inst_ack_0, ack => testConfigure_CP_0_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	341 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	50 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_125_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_125_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_125_Update/ca
      -- 
    ca_331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_125_inst_ack_1, ack => testConfigure_CP_0_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	341 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	50 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_final_index_sum_regn_sample_complete
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_final_index_sum_regn_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_final_index_sum_regn_Sample/ack
      -- 
    ack_357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_131_index_offset_ack_0, ack => testConfigure_CP_0_elements(26)); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	341 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (11) 
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_root_address_calculated
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_offset_calculated
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/addr_of_132_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_final_index_sum_regn_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_final_index_sum_regn_Update/ack
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_base_plus_offset/$entry
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_base_plus_offset/$exit
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_base_plus_offset/sum_rename_req
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_base_plus_offset/sum_rename_ack
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/addr_of_132_request/$entry
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/addr_of_132_request/req
      -- 
    ack_362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_131_index_offset_ack_1, ack => testConfigure_CP_0_elements(27)); -- 
    req_371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(27), ack => addr_of_132_final_reg_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/addr_of_132_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/addr_of_132_request/$exit
      -- CP-element group 28: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/addr_of_132_request/ack
      -- 
    ack_372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_132_final_reg_ack_0, ack => testConfigure_CP_0_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	341 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: 	36 
    -- CP-element group 29:  members (44) 
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/addr_of_132_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/addr_of_132_complete/$exit
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/addr_of_132_complete/ack
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_base_address_calculated
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_word_address_calculated
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_root_address_calculated
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_base_address_resized
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_base_addr_resize/$entry
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_base_addr_resize/$exit
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_base_addr_resize/base_resize_req
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_base_addr_resize/base_resize_ack
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_base_plus_offset/$entry
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_base_plus_offset/$exit
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_base_plus_offset/sum_rename_req
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_base_plus_offset/sum_rename_ack
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_word_addrgen/$entry
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_word_addrgen/$exit
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_word_addrgen/root_register_req
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_word_addrgen/root_register_ack
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_Sample/ptr_deref_135_Split/$entry
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_Sample/ptr_deref_135_Split/$exit
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_Sample/ptr_deref_135_Split/split_req
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_Sample/ptr_deref_135_Split/split_ack
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_Sample/word_access_start/$entry
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_Sample/word_access_start/word_0/$entry
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_Sample/word_access_start/word_0/rr
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_base_address_calculated
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_word_address_calculated
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_root_address_calculated
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_base_address_resized
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_base_addr_resize/$entry
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_base_addr_resize/$exit
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_base_addr_resize/base_resize_req
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_base_addr_resize/base_resize_ack
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_base_plus_offset/$entry
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_base_plus_offset/$exit
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_base_plus_offset/sum_rename_req
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_base_plus_offset/sum_rename_ack
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_word_addrgen/$entry
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_word_addrgen/$exit
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_word_addrgen/root_register_req
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_word_addrgen/root_register_ack
      -- 
    ack_377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_132_final_reg_ack_1, ack => testConfigure_CP_0_elements(29)); -- 
    rr_415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(29), ack => ptr_deref_135_store_0_req_0); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	48 
    -- CP-element group 30:  members (5) 
      -- CP-element group 30: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_Sample/word_access_start/$exit
      -- CP-element group 30: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_Sample/word_access_start/word_0/$exit
      -- CP-element group 30: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_Sample/word_access_start/word_0/ra
      -- 
    ra_416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_135_store_0_ack_0, ack => testConfigure_CP_0_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	341 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	50 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_Update/word_access_complete/$exit
      -- CP-element group 31: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_Update/word_access_complete/word_0/$exit
      -- CP-element group 31: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_Update/word_access_complete/word_0/ca
      -- 
    ca_427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_135_store_0_ack_1, ack => testConfigure_CP_0_elements(31)); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	341 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_145_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_145_update_start_
      -- CP-element group 32: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_145_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_145_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_145_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_145_Update/cr
      -- 
    ra_436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_145_inst_ack_0, ack => testConfigure_CP_0_elements(32)); -- 
    cr_440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(32), ack => RPIPE_ConvTranspose_input_pipe_145_inst_req_1); -- 
    -- CP-element group 33:  fork  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	44 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (9) 
      -- CP-element group 33: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_145_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_145_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_145_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_149_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_149_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_149_Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_189_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_189_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_189_Sample/rr
      -- 
    ca_441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_145_inst_ack_1, ack => testConfigure_CP_0_elements(33)); -- 
    rr_577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(33), ack => RPIPE_ConvTranspose_input_pipe_189_inst_req_0); -- 
    rr_449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(33), ack => type_cast_149_inst_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_149_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_149_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_149_Sample/ra
      -- 
    ra_450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_149_inst_ack_0, ack => testConfigure_CP_0_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	341 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_149_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_149_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_149_Update/ca
      -- 
    ca_455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_149_inst_ack_1, ack => testConfigure_CP_0_elements(35)); -- 
    -- CP-element group 36:  join  transition  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	29 
    -- CP-element group 36: 	35 
    -- CP-element group 36: 	48 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (9) 
      -- CP-element group 36: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_Sample/ptr_deref_157_Split/$entry
      -- CP-element group 36: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_Sample/ptr_deref_157_Split/$exit
      -- CP-element group 36: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_Sample/ptr_deref_157_Split/split_req
      -- CP-element group 36: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_Sample/ptr_deref_157_Split/split_ack
      -- CP-element group 36: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_Sample/word_access_start/$entry
      -- CP-element group 36: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_Sample/word_access_start/word_0/$entry
      -- CP-element group 36: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_Sample/word_access_start/word_0/rr
      -- 
    rr_493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(36), ack => ptr_deref_157_store_0_req_0); -- 
    testConfigure_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(29) & testConfigure_CP_0_elements(35) & testConfigure_CP_0_elements(48);
      gj_testConfigure_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	49 
    -- CP-element group 37:  members (5) 
      -- CP-element group 37: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_Sample/word_access_start/$exit
      -- CP-element group 37: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_Sample/word_access_start/word_0/$exit
      -- CP-element group 37: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_Sample/word_access_start/word_0/ra
      -- 
    ra_494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_157_store_0_ack_0, ack => testConfigure_CP_0_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	341 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	50 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_Update/word_access_complete/$exit
      -- CP-element group 38: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_Update/word_access_complete/word_0/$exit
      -- CP-element group 38: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_Update/word_access_complete/word_0/ca
      -- 
    ca_505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_157_store_0_ack_1, ack => testConfigure_CP_0_elements(38)); -- 
    -- CP-element group 39:  join  transition  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	49 
    -- CP-element group 39: 	341 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (5) 
      -- CP-element group 39: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_Sample/word_access_start/$entry
      -- CP-element group 39: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_Sample/word_access_start/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_Sample/word_access_start/word_0/rr
      -- 
    rr_538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(39), ack => ptr_deref_174_load_0_req_0); -- 
    testConfigure_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(49) & testConfigure_CP_0_elements(341);
      gj_testConfigure_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_Sample/word_access_start/$exit
      -- CP-element group 40: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_Sample/word_access_start/word_0/$exit
      -- CP-element group 40: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_Sample/word_access_start/word_0/ra
      -- 
    ra_539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_174_load_0_ack_0, ack => testConfigure_CP_0_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	341 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (12) 
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_Update/word_access_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_Update/word_access_complete/word_0/$exit
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_Update/word_access_complete/word_0/ca
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_Update/ptr_deref_174_Merge/$entry
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_Update/ptr_deref_174_Merge/$exit
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_Update/ptr_deref_174_Merge/merge_req
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_Update/ptr_deref_174_Merge/merge_ack
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_178_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_178_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_178_Sample/rr
      -- 
    ca_550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_174_load_0_ack_1, ack => testConfigure_CP_0_elements(41)); -- 
    rr_563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(41), ack => type_cast_178_inst_req_0); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_178_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_178_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_178_Sample/ra
      -- 
    ra_564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_178_inst_ack_0, ack => testConfigure_CP_0_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	341 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	50 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_178_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_178_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_178_Update/ca
      -- 
    ca_569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_178_inst_ack_1, ack => testConfigure_CP_0_elements(43)); -- 
    -- CP-element group 44:  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	33 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (6) 
      -- CP-element group 44: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_189_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_189_update_start_
      -- CP-element group 44: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_189_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_189_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_189_Update/$entry
      -- CP-element group 44: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_189_Update/cr
      -- 
    ra_578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_189_inst_ack_0, ack => testConfigure_CP_0_elements(44)); -- 
    cr_582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(44), ack => RPIPE_ConvTranspose_input_pipe_189_inst_req_1); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_189_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_189_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_189_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_193_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_193_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_193_Sample/rr
      -- 
    ca_583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_189_inst_ack_1, ack => testConfigure_CP_0_elements(45)); -- 
    rr_591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(45), ack => type_cast_193_inst_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_193_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_193_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_193_Sample/ra
      -- 
    ra_592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_193_inst_ack_0, ack => testConfigure_CP_0_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	341 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	50 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_193_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_193_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_193_Update/ca
      -- 
    ca_597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_193_inst_ack_1, ack => testConfigure_CP_0_elements(47)); -- 
    -- CP-element group 48:  transition  delay-element  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	30 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	36 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_ptr_deref_157_delay
      -- 
    -- Element group testConfigure_CP_0_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(30), ack => testConfigure_CP_0_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  transition  delay-element  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	37 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	39 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_ptr_deref_174_delay
      -- 
    -- Element group testConfigure_CP_0_elements(49) is a control-delay.
    cp_element_49_delay: control_delay_element  generic map(name => " 49_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(37), ack => testConfigure_CP_0_elements(49), clk => clk, reset =>reset);
    -- CP-element group 50:  branch  join  transition  place  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	43 
    -- CP-element group 50: 	25 
    -- CP-element group 50: 	26 
    -- CP-element group 50: 	31 
    -- CP-element group 50: 	38 
    -- CP-element group 50: 	47 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (10) 
      -- CP-element group 50: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194__exit__
      -- CP-element group 50: 	 branch_block_stmt_34/if_stmt_195__entry__
      -- CP-element group 50: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/$exit
      -- CP-element group 50: 	 branch_block_stmt_34/if_stmt_195_dead_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_34/if_stmt_195_eval_test/$entry
      -- CP-element group 50: 	 branch_block_stmt_34/if_stmt_195_eval_test/$exit
      -- CP-element group 50: 	 branch_block_stmt_34/if_stmt_195_eval_test/branch_req
      -- CP-element group 50: 	 branch_block_stmt_34/R_cmp_196_place
      -- CP-element group 50: 	 branch_block_stmt_34/if_stmt_195_if_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_34/if_stmt_195_else_link/$entry
      -- 
    branch_req_607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(50), ack => if_stmt_195_branch_req_0); -- 
    testConfigure_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(43) & testConfigure_CP_0_elements(25) & testConfigure_CP_0_elements(26) & testConfigure_CP_0_elements(31) & testConfigure_CP_0_elements(38) & testConfigure_CP_0_elements(47);
      gj_testConfigure_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  fork  transition  place  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	326 
    -- CP-element group 51: 	327 
    -- CP-element group 51: 	329 
    -- CP-element group 51: 	330 
    -- CP-element group 51:  members (20) 
      -- CP-element group 51: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_115/SplitProtocol/Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_34/if_stmt_195_if_link/$exit
      -- CP-element group 51: 	 branch_block_stmt_34/if_stmt_195_if_link/if_choice_transition
      -- CP-element group 51: 	 branch_block_stmt_34/forx_xbody_forx_xbody
      -- CP-element group 51: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_115/SplitProtocol/Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_115/SplitProtocol/Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_115/SplitProtocol/$entry
      -- CP-element group 51: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_115/$entry
      -- CP-element group 51: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/$entry
      -- CP-element group 51: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_110/$entry
      -- CP-element group 51: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_115/SplitProtocol/Update/cr
      -- CP-element group 51: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_103/phi_stmt_103_sources/type_cast_106/SplitProtocol/Update/cr
      -- CP-element group 51: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_103/phi_stmt_103_sources/type_cast_106/SplitProtocol/Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_103/phi_stmt_103_sources/type_cast_106/SplitProtocol/Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_103/phi_stmt_103_sources/type_cast_106/SplitProtocol/Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_103/phi_stmt_103_sources/type_cast_106/SplitProtocol/$entry
      -- CP-element group 51: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_103/phi_stmt_103_sources/type_cast_106/$entry
      -- CP-element group 51: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_103/phi_stmt_103_sources/$entry
      -- CP-element group 51: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_103/$entry
      -- CP-element group 51: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/$entry
      -- 
    if_choice_transition_612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_195_branch_ack_1, ack => testConfigure_CP_0_elements(51)); -- 
    rr_3520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(51), ack => type_cast_115_inst_req_0); -- 
    cr_3525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(51), ack => type_cast_115_inst_req_1); -- 
    cr_3502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(51), ack => type_cast_106_inst_req_1); -- 
    rr_3497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(51), ack => type_cast_106_inst_req_0); -- 
    -- CP-element group 52:  fork  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	342 
    -- CP-element group 52: 	343 
    -- CP-element group 52:  members (12) 
      -- CP-element group 52: 	 branch_block_stmt_34/if_stmt_195_else_link/$exit
      -- CP-element group 52: 	 branch_block_stmt_34/if_stmt_195_else_link/else_choice_transition
      -- CP-element group 52: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 52: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_202/phi_stmt_202_sources/type_cast_205/SplitProtocol/$entry
      -- CP-element group 52: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_202/phi_stmt_202_sources/type_cast_205/SplitProtocol/Update/cr
      -- CP-element group 52: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_202/phi_stmt_202_sources/type_cast_205/SplitProtocol/Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_202/phi_stmt_202_sources/type_cast_205/SplitProtocol/Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_202/phi_stmt_202_sources/type_cast_205/SplitProtocol/Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_202/phi_stmt_202_sources/type_cast_205/$entry
      -- CP-element group 52: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_202/phi_stmt_202_sources/$entry
      -- CP-element group 52: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_202/$entry
      -- CP-element group 52: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- 
    else_choice_transition_616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_195_branch_ack_0, ack => testConfigure_CP_0_elements(52)); -- 
    cr_3595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(52), ack => type_cast_205_inst_req_1); -- 
    rr_3590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(52), ack => type_cast_205_inst_req_0); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	353 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	62 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_Sample/word_access_start/$exit
      -- CP-element group 53: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_Sample/word_access_start/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_Sample/word_access_start/word_0/ra
      -- 
    ra_660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_223_store_0_ack_0, ack => testConfigure_CP_0_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	353 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	63 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_Update/word_access_complete/$exit
      -- CP-element group 54: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_Update/word_access_complete/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_Update/word_access_complete/word_0/ca
      -- 
    ca_671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_223_store_0_ack_1, ack => testConfigure_CP_0_elements(54)); -- 
    -- CP-element group 55:  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	353 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (6) 
      -- CP-element group 55: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/RPIPE_ConvTranspose_input_pipe_233_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/RPIPE_ConvTranspose_input_pipe_233_update_start_
      -- CP-element group 55: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/RPIPE_ConvTranspose_input_pipe_233_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/RPIPE_ConvTranspose_input_pipe_233_Sample/ra
      -- CP-element group 55: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/RPIPE_ConvTranspose_input_pipe_233_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/RPIPE_ConvTranspose_input_pipe_233_Update/cr
      -- 
    ra_680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_233_inst_ack_0, ack => testConfigure_CP_0_elements(55)); -- 
    cr_684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(55), ack => RPIPE_ConvTranspose_input_pipe_233_inst_req_1); -- 
    -- CP-element group 56:  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (6) 
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/RPIPE_ConvTranspose_input_pipe_233_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/RPIPE_ConvTranspose_input_pipe_233_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/RPIPE_ConvTranspose_input_pipe_233_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/type_cast_237_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/type_cast_237_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/type_cast_237_Sample/rr
      -- 
    ca_685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_233_inst_ack_1, ack => testConfigure_CP_0_elements(56)); -- 
    rr_693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => type_cast_237_inst_req_0); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/type_cast_237_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/type_cast_237_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/type_cast_237_Sample/ra
      -- 
    ra_694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_237_inst_ack_0, ack => testConfigure_CP_0_elements(57)); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	353 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/type_cast_237_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/type_cast_237_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/type_cast_237_Update/ca
      -- 
    ca_699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_237_inst_ack_1, ack => testConfigure_CP_0_elements(58)); -- 
    -- CP-element group 59:  join  transition  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: 	62 
    -- CP-element group 59: 	353 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (9) 
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_Sample/ptr_deref_251_Split/$entry
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_Sample/ptr_deref_251_Split/$exit
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_Sample/ptr_deref_251_Split/split_req
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_Sample/ptr_deref_251_Split/split_ack
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_Sample/word_access_start/$entry
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_Sample/word_access_start/word_0/$entry
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_Sample/word_access_start/word_0/rr
      -- 
    rr_737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(59), ack => ptr_deref_251_store_0_req_0); -- 
    testConfigure_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(58) & testConfigure_CP_0_elements(62) & testConfigure_CP_0_elements(353);
      gj_testConfigure_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (5) 
      -- CP-element group 60: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_Sample/word_access_start/$exit
      -- CP-element group 60: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_Sample/word_access_start/word_0/$exit
      -- CP-element group 60: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_Sample/word_access_start/word_0/ra
      -- 
    ra_738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_251_store_0_ack_0, ack => testConfigure_CP_0_elements(60)); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	353 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (5) 
      -- CP-element group 61: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_Update/word_access_complete/$exit
      -- CP-element group 61: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_Update/word_access_complete/word_0/$exit
      -- CP-element group 61: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_Update/word_access_complete/word_0/ca
      -- 
    ca_749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_251_store_0_ack_1, ack => testConfigure_CP_0_elements(61)); -- 
    -- CP-element group 62:  transition  delay-element  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	53 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	59 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_ptr_deref_251_delay
      -- 
    -- Element group testConfigure_CP_0_elements(62) is a control-delay.
    cp_element_62_delay: control_delay_element  generic map(name => " 62_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(53), ack => testConfigure_CP_0_elements(62), clk => clk, reset =>reset);
    -- CP-element group 63:  branch  join  transition  place  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	54 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (10) 
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259__exit__
      -- CP-element group 63: 	 branch_block_stmt_34/if_stmt_260__entry__
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/$exit
      -- CP-element group 63: 	 branch_block_stmt_34/if_stmt_260_dead_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_34/if_stmt_260_eval_test/$entry
      -- CP-element group 63: 	 branch_block_stmt_34/if_stmt_260_eval_test/$exit
      -- CP-element group 63: 	 branch_block_stmt_34/if_stmt_260_eval_test/branch_req
      -- CP-element group 63: 	 branch_block_stmt_34/R_cmp40311_261_place
      -- CP-element group 63: 	 branch_block_stmt_34/if_stmt_260_if_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_34/if_stmt_260_else_link/$entry
      -- 
    branch_req_758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(63), ack => if_stmt_260_branch_req_0); -- 
    testConfigure_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(54) & testConfigure_CP_0_elements(61);
      gj_testConfigure_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  place  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	360 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_34/if_stmt_260_if_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_34/if_stmt_260_if_link/if_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_34/forx_xend_bbx_xnph307
      -- CP-element group 64: 	 branch_block_stmt_34/forx_xend_bbx_xnph307_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_34/forx_xend_bbx_xnph307_PhiReq/$exit
      -- 
    if_choice_transition_763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_260_branch_ack_1, ack => testConfigure_CP_0_elements(64)); -- 
    -- CP-element group 65:  merge  transition  place  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	357 
    -- CP-element group 65:  members (14) 
      -- CP-element group 65: 	 branch_block_stmt_34/merge_stmt_266__exit__
      -- CP-element group 65: 	 branch_block_stmt_34/forx_xbody42x_xpreheader_forx_xbody42
      -- CP-element group 65: 	 branch_block_stmt_34/if_stmt_260_else_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_34/if_stmt_260_else_link/else_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_34/forx_xend_forx_xbody42x_xpreheader
      -- CP-element group 65: 	 branch_block_stmt_34/forx_xend_forx_xbody42x_xpreheader_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_34/forx_xend_forx_xbody42x_xpreheader_PhiReq/$exit
      -- CP-element group 65: 	 branch_block_stmt_34/merge_stmt_266_PhiReqMerge
      -- CP-element group 65: 	 branch_block_stmt_34/merge_stmt_266_PhiAck/$entry
      -- CP-element group 65: 	 branch_block_stmt_34/merge_stmt_266_PhiAck/$exit
      -- CP-element group 65: 	 branch_block_stmt_34/merge_stmt_266_PhiAck/dummy
      -- CP-element group 65: 	 branch_block_stmt_34/forx_xbody42x_xpreheader_forx_xbody42_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_34/forx_xbody42x_xpreheader_forx_xbody42_PhiReq/phi_stmt_269/$entry
      -- CP-element group 65: 	 branch_block_stmt_34/forx_xbody42x_xpreheader_forx_xbody42_PhiReq/phi_stmt_269/phi_stmt_269_sources/$entry
      -- 
    else_choice_transition_767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_260_branch_ack_0, ack => testConfigure_CP_0_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	359 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_285_Sample/ra
      -- CP-element group 66: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_285_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_285_Sample/$exit
      -- 
    ra_781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_285_inst_ack_0, ack => testConfigure_CP_0_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	359 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	93 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_285_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_285_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_285_update_completed_
      -- 
    ca_786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_285_inst_ack_1, ack => testConfigure_CP_0_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	359 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	93 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_final_index_sum_regn_sample_complete
      -- CP-element group 68: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_final_index_sum_regn_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_final_index_sum_regn_Sample/ack
      -- 
    ack_812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_291_index_offset_ack_0, ack => testConfigure_CP_0_elements(68)); -- 
    -- CP-element group 69:  transition  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	359 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (11) 
      -- CP-element group 69: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/addr_of_292_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_root_address_calculated
      -- CP-element group 69: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_offset_calculated
      -- CP-element group 69: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_final_index_sum_regn_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_final_index_sum_regn_Update/ack
      -- CP-element group 69: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_base_plus_offset/$entry
      -- CP-element group 69: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_base_plus_offset/$exit
      -- CP-element group 69: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_base_plus_offset/sum_rename_req
      -- CP-element group 69: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_base_plus_offset/sum_rename_ack
      -- CP-element group 69: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/addr_of_292_request/$entry
      -- CP-element group 69: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/addr_of_292_request/req
      -- 
    ack_817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_291_index_offset_ack_1, ack => testConfigure_CP_0_elements(69)); -- 
    req_826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(69), ack => addr_of_292_final_reg_req_0); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/addr_of_292_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/addr_of_292_request/$exit
      -- CP-element group 70: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/addr_of_292_request/ack
      -- 
    ack_827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_292_final_reg_ack_0, ack => testConfigure_CP_0_elements(70)); -- 
    -- CP-element group 71:  fork  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	359 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	76 
    -- CP-element group 71: 	83 
    -- CP-element group 71:  members (35) 
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/addr_of_292_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/addr_of_292_complete/$exit
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/addr_of_292_complete/ack
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_base_address_calculated
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_word_address_calculated
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_root_address_calculated
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_base_address_resized
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_base_addr_resize/$entry
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_base_addr_resize/$exit
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_base_addr_resize/base_resize_req
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_base_addr_resize/base_resize_ack
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_base_plus_offset/$entry
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_base_plus_offset/$exit
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_base_plus_offset/sum_rename_req
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_base_plus_offset/sum_rename_ack
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_word_addrgen/$entry
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_word_addrgen/$exit
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_word_addrgen/root_register_req
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_word_addrgen/root_register_ack
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_base_address_calculated
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_word_address_calculated
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_root_address_calculated
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_base_address_resized
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_base_addr_resize/$entry
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_base_addr_resize/$exit
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_base_addr_resize/base_resize_req
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_base_addr_resize/base_resize_ack
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_base_plus_offset/$entry
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_base_plus_offset/$exit
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_base_plus_offset/sum_rename_req
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_base_plus_offset/sum_rename_ack
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_word_addrgen/$entry
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_word_addrgen/$exit
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_word_addrgen/root_register_req
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_word_addrgen/root_register_ack
      -- 
    ack_832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_292_final_reg_ack_1, ack => testConfigure_CP_0_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	359 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_295_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_295_update_start_
      -- CP-element group 72: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_295_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_295_Sample/ra
      -- CP-element group 72: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_295_Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_295_Update/cr
      -- 
    ra_841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_295_inst_ack_0, ack => testConfigure_CP_0_elements(72)); -- 
    cr_845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(72), ack => RPIPE_ConvTranspose_input_pipe_295_inst_req_1); -- 
    -- CP-element group 73:  fork  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73: 	79 
    -- CP-element group 73:  members (9) 
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_295_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_295_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_295_Update/ca
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_299_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_299_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_299_Sample/rr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_312_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_312_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_312_Sample/rr
      -- 
    ca_846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_295_inst_ack_1, ack => testConfigure_CP_0_elements(73)); -- 
    rr_854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => type_cast_299_inst_req_0); -- 
    rr_918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => RPIPE_ConvTranspose_input_pipe_312_inst_req_0); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_299_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_299_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_299_Sample/ra
      -- 
    ra_855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_299_inst_ack_0, ack => testConfigure_CP_0_elements(74)); -- 
    -- CP-element group 75:  fork  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	359 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75: 	83 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_299_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_299_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_299_Update/ca
      -- 
    ca_860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_299_inst_ack_1, ack => testConfigure_CP_0_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	71 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (9) 
      -- CP-element group 76: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_Sample/ptr_deref_302_Split/$entry
      -- CP-element group 76: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_Sample/ptr_deref_302_Split/$exit
      -- CP-element group 76: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_Sample/ptr_deref_302_Split/split_req
      -- CP-element group 76: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_Sample/ptr_deref_302_Split/split_ack
      -- CP-element group 76: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_Sample/word_access_start/$entry
      -- CP-element group 76: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_Sample/word_access_start/word_0/$entry
      -- CP-element group 76: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_Sample/word_access_start/word_0/rr
      -- 
    rr_898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(76), ack => ptr_deref_302_store_0_req_0); -- 
    testConfigure_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(71) & testConfigure_CP_0_elements(75);
      gj_testConfigure_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	91 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_Sample/word_access_start/$exit
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_Sample/word_access_start/word_0/$exit
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_Sample/word_access_start/word_0/ra
      -- 
    ra_899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_302_store_0_ack_0, ack => testConfigure_CP_0_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	359 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	93 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_Update/word_access_complete/$exit
      -- CP-element group 78: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_Update/word_access_complete/word_0/$exit
      -- CP-element group 78: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_Update/word_access_complete/word_0/ca
      -- 
    ca_910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_302_store_0_ack_1, ack => testConfigure_CP_0_elements(78)); -- 
    -- CP-element group 79:  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	73 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (6) 
      -- CP-element group 79: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_312_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_312_update_start_
      -- CP-element group 79: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_312_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_312_Sample/ra
      -- CP-element group 79: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_312_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_312_Update/cr
      -- 
    ra_919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_312_inst_ack_0, ack => testConfigure_CP_0_elements(79)); -- 
    cr_923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(79), ack => RPIPE_ConvTranspose_input_pipe_312_inst_req_1); -- 
    -- CP-element group 80:  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (6) 
      -- CP-element group 80: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_312_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_312_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_312_Update/ca
      -- CP-element group 80: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_316_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_316_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_316_Sample/rr
      -- 
    ca_924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_312_inst_ack_1, ack => testConfigure_CP_0_elements(80)); -- 
    rr_932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(80), ack => type_cast_316_inst_req_0); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_316_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_316_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_316_Sample/ra
      -- 
    ra_933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_316_inst_ack_0, ack => testConfigure_CP_0_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	359 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_316_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_316_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_316_Update/ca
      -- 
    ca_938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_316_inst_ack_1, ack => testConfigure_CP_0_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	71 
    -- CP-element group 83: 	75 
    -- CP-element group 83: 	82 
    -- CP-element group 83: 	91 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_Sample/ptr_deref_324_Split/$entry
      -- CP-element group 83: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_Sample/ptr_deref_324_Split/$exit
      -- CP-element group 83: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_Sample/ptr_deref_324_Split/split_req
      -- CP-element group 83: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_Sample/ptr_deref_324_Split/split_ack
      -- CP-element group 83: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_Sample/word_access_start/$entry
      -- CP-element group 83: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_Sample/word_access_start/word_0/$entry
      -- CP-element group 83: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_Sample/word_access_start/word_0/rr
      -- 
    rr_976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(83), ack => ptr_deref_324_store_0_req_0); -- 
    testConfigure_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(71) & testConfigure_CP_0_elements(75) & testConfigure_CP_0_elements(82) & testConfigure_CP_0_elements(91);
      gj_testConfigure_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	92 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_Sample/word_access_start/$exit
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_Sample/word_access_start/word_0/$exit
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_Sample/word_access_start/word_0/ra
      -- 
    ra_977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_324_store_0_ack_0, ack => testConfigure_CP_0_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	359 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	93 
    -- CP-element group 85:  members (5) 
      -- CP-element group 85: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_Update/word_access_complete/$exit
      -- CP-element group 85: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_Update/word_access_complete/word_0/$exit
      -- CP-element group 85: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_Update/word_access_complete/word_0/ca
      -- 
    ca_988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_324_store_0_ack_1, ack => testConfigure_CP_0_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	92 
    -- CP-element group 86: 	359 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_Sample/word_access_start/$entry
      -- CP-element group 86: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_Sample/word_access_start/word_0/$entry
      -- CP-element group 86: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_Sample/word_access_start/word_0/rr
      -- 
    rr_1021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(86), ack => ptr_deref_341_load_0_req_0); -- 
    testConfigure_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(92) & testConfigure_CP_0_elements(359);
      gj_testConfigure_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_Sample/word_access_start/$exit
      -- CP-element group 87: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_Sample/word_access_start/word_0/$exit
      -- CP-element group 87: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_Sample/word_access_start/word_0/ra
      -- 
    ra_1022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_341_load_0_ack_0, ack => testConfigure_CP_0_elements(87)); -- 
    -- CP-element group 88:  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	359 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (12) 
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_Update/word_access_complete/$exit
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_Update/word_access_complete/word_0/$exit
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_Update/word_access_complete/word_0/ca
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_Update/ptr_deref_341_Merge/$entry
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_Update/ptr_deref_341_Merge/$exit
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_Update/ptr_deref_341_Merge/merge_req
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_Update/ptr_deref_341_Merge/merge_ack
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_345_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_345_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_345_Sample/rr
      -- 
    ca_1033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_341_load_0_ack_1, ack => testConfigure_CP_0_elements(88)); -- 
    rr_1046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(88), ack => type_cast_345_inst_req_0); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_345_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_345_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_345_Sample/ra
      -- 
    ra_1047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_345_inst_ack_0, ack => testConfigure_CP_0_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	359 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	93 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_345_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_345_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_345_Update/ca
      -- 
    ca_1052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_345_inst_ack_1, ack => testConfigure_CP_0_elements(90)); -- 
    -- CP-element group 91:  transition  delay-element  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	77 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	83 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_ptr_deref_324_delay
      -- 
    -- Element group testConfigure_CP_0_elements(91) is a control-delay.
    cp_element_91_delay: control_delay_element  generic map(name => " 91_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(77), ack => testConfigure_CP_0_elements(91), clk => clk, reset =>reset);
    -- CP-element group 92:  transition  delay-element  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	84 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	86 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_ptr_deref_341_delay
      -- 
    -- Element group testConfigure_CP_0_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(84), ack => testConfigure_CP_0_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  branch  join  transition  place  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	67 
    -- CP-element group 93: 	68 
    -- CP-element group 93: 	78 
    -- CP-element group 93: 	85 
    -- CP-element group 93: 	90 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (10) 
      -- CP-element group 93: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353__exit__
      -- CP-element group 93: 	 branch_block_stmt_34/if_stmt_354__entry__
      -- CP-element group 93: 	 branch_block_stmt_34/if_stmt_354_else_link/$entry
      -- CP-element group 93: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/$exit
      -- CP-element group 93: 	 branch_block_stmt_34/R_cmp40_355_place
      -- CP-element group 93: 	 branch_block_stmt_34/if_stmt_354_if_link/$entry
      -- CP-element group 93: 	 branch_block_stmt_34/if_stmt_354_dead_link/$entry
      -- CP-element group 93: 	 branch_block_stmt_34/if_stmt_354_eval_test/$entry
      -- CP-element group 93: 	 branch_block_stmt_34/if_stmt_354_eval_test/$exit
      -- CP-element group 93: 	 branch_block_stmt_34/if_stmt_354_eval_test/branch_req
      -- 
    branch_req_1062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(93), ack => if_stmt_354_branch_req_0); -- 
    testConfigure_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(67) & testConfigure_CP_0_elements(68) & testConfigure_CP_0_elements(78) & testConfigure_CP_0_elements(85) & testConfigure_CP_0_elements(90);
      gj_testConfigure_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  fork  transition  place  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	354 
    -- CP-element group 94: 	355 
    -- CP-element group 94:  members (12) 
      -- CP-element group 94: 	 branch_block_stmt_34/if_stmt_354_if_link/$exit
      -- CP-element group 94: 	 branch_block_stmt_34/if_stmt_354_if_link/if_choice_transition
      -- CP-element group 94: 	 branch_block_stmt_34/forx_xbody42_forx_xbody42
      -- CP-element group 94: 	 branch_block_stmt_34/forx_xbody42_forx_xbody42_PhiReq/$entry
      -- CP-element group 94: 	 branch_block_stmt_34/forx_xbody42_forx_xbody42_PhiReq/phi_stmt_269/$entry
      -- CP-element group 94: 	 branch_block_stmt_34/forx_xbody42_forx_xbody42_PhiReq/phi_stmt_269/phi_stmt_269_sources/$entry
      -- CP-element group 94: 	 branch_block_stmt_34/forx_xbody42_forx_xbody42_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_272/$entry
      -- CP-element group 94: 	 branch_block_stmt_34/forx_xbody42_forx_xbody42_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_272/SplitProtocol/$entry
      -- CP-element group 94: 	 branch_block_stmt_34/forx_xbody42_forx_xbody42_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_272/SplitProtocol/Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_34/forx_xbody42_forx_xbody42_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_272/SplitProtocol/Sample/rr
      -- CP-element group 94: 	 branch_block_stmt_34/forx_xbody42_forx_xbody42_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_272/SplitProtocol/Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_34/forx_xbody42_forx_xbody42_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_272/SplitProtocol/Update/cr
      -- 
    if_choice_transition_1067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_354_branch_ack_1, ack => testConfigure_CP_0_elements(94)); -- 
    rr_3690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(94), ack => type_cast_272_inst_req_0); -- 
    cr_3695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(94), ack => type_cast_272_inst_req_1); -- 
    -- CP-element group 95:  merge  transition  place  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	360 
    -- CP-element group 95:  members (13) 
      -- CP-element group 95: 	 branch_block_stmt_34/merge_stmt_360__exit__
      -- CP-element group 95: 	 branch_block_stmt_34/bbx_xnph307x_xloopexit_bbx_xnph307
      -- CP-element group 95: 	 branch_block_stmt_34/forx_xbody42_bbx_xnph307x_xloopexit
      -- CP-element group 95: 	 branch_block_stmt_34/if_stmt_354_else_link/else_choice_transition
      -- CP-element group 95: 	 branch_block_stmt_34/if_stmt_354_else_link/$exit
      -- CP-element group 95: 	 branch_block_stmt_34/forx_xbody42_bbx_xnph307x_xloopexit_PhiReq/$entry
      -- CP-element group 95: 	 branch_block_stmt_34/forx_xbody42_bbx_xnph307x_xloopexit_PhiReq/$exit
      -- CP-element group 95: 	 branch_block_stmt_34/merge_stmt_360_PhiReqMerge
      -- CP-element group 95: 	 branch_block_stmt_34/merge_stmt_360_PhiAck/$entry
      -- CP-element group 95: 	 branch_block_stmt_34/merge_stmt_360_PhiAck/$exit
      -- CP-element group 95: 	 branch_block_stmt_34/merge_stmt_360_PhiAck/dummy
      -- CP-element group 95: 	 branch_block_stmt_34/bbx_xnph307x_xloopexit_bbx_xnph307_PhiReq/$entry
      -- CP-element group 95: 	 branch_block_stmt_34/bbx_xnph307x_xloopexit_bbx_xnph307_PhiReq/$exit
      -- 
    else_choice_transition_1071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_354_branch_ack_0, ack => testConfigure_CP_0_elements(95)); -- 
    -- CP-element group 96:  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	360 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (6) 
      -- CP-element group 96: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/RPIPE_ConvTranspose_input_pipe_364_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/RPIPE_ConvTranspose_input_pipe_364_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/RPIPE_ConvTranspose_input_pipe_364_update_start_
      -- CP-element group 96: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/RPIPE_ConvTranspose_input_pipe_364_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/RPIPE_ConvTranspose_input_pipe_364_Update/cr
      -- CP-element group 96: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/RPIPE_ConvTranspose_input_pipe_364_Update/$entry
      -- 
    ra_1085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_364_inst_ack_0, ack => testConfigure_CP_0_elements(96)); -- 
    cr_1089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(96), ack => RPIPE_ConvTranspose_input_pipe_364_inst_req_1); -- 
    -- CP-element group 97:  transition  input  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (6) 
      -- CP-element group 97: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/RPIPE_ConvTranspose_input_pipe_364_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/type_cast_368_Sample/rr
      -- CP-element group 97: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/type_cast_368_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/type_cast_368_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/RPIPE_ConvTranspose_input_pipe_364_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/RPIPE_ConvTranspose_input_pipe_364_Update/$exit
      -- 
    ca_1090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_364_inst_ack_1, ack => testConfigure_CP_0_elements(97)); -- 
    rr_1098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(97), ack => type_cast_368_inst_req_0); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/type_cast_368_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/type_cast_368_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/type_cast_368_sample_completed_
      -- 
    ra_1099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_368_inst_ack_0, ack => testConfigure_CP_0_elements(98)); -- 
    -- CP-element group 99:  fork  transition  place  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	360 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	361 
    -- CP-element group 99: 	362 
    -- CP-element group 99: 	363 
    -- CP-element group 99:  members (17) 
      -- CP-element group 99: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369__exit__
      -- CP-element group 99: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69
      -- CP-element group 99: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/type_cast_368_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/type_cast_368_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/type_cast_368_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/$exit
      -- CP-element group 99: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/$entry
      -- CP-element group 99: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_372/$entry
      -- CP-element group 99: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_372/phi_stmt_372_sources/$entry
      -- CP-element group 99: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_379/$entry
      -- CP-element group 99: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/$entry
      -- CP-element group 99: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_382/$entry
      -- CP-element group 99: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_382/SplitProtocol/$entry
      -- CP-element group 99: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_382/SplitProtocol/Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_382/SplitProtocol/Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_382/SplitProtocol/Update/$entry
      -- CP-element group 99: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_382/SplitProtocol/Update/cr
      -- 
    ca_1104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_368_inst_ack_1, ack => testConfigure_CP_0_elements(99)); -- 
    rr_3763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(99), ack => type_cast_382_inst_req_0); -- 
    cr_3768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(99), ack => type_cast_382_inst_req_1); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	376 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/addr_of_389_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/addr_of_389_request/ack
      -- CP-element group 100: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/addr_of_389_request/$exit
      -- 
    ack_1141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_389_final_reg_ack_0, ack => testConfigure_CP_0_elements(100)); -- 
    -- CP-element group 101:  join  fork  transition  input  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	376 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101: 	108 
    -- CP-element group 101:  members (44) 
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_word_addrgen/root_register_ack
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_base_address_resized
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_root_address_calculated
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_word_address_calculated
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_sample_start_
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/addr_of_389_complete/ack
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/addr_of_389_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_Sample/word_access_start/word_0/rr
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_Sample/word_access_start/word_0/$entry
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_base_address_calculated
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_Sample/word_access_start/$entry
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_word_addrgen/root_register_req
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_Sample/ptr_deref_392_Split/split_ack
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_Sample/ptr_deref_392_Split/split_req
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_Sample/ptr_deref_392_Split/$exit
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_word_addrgen/$exit
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_Sample/ptr_deref_392_Split/$entry
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/addr_of_389_complete/$exit
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_word_addrgen/$entry
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_base_plus_offset/sum_rename_ack
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_word_addrgen/root_register_ack
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_base_plus_offset/sum_rename_req
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_word_addrgen/root_register_req
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_word_addrgen/$exit
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_word_addrgen/$entry
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_base_plus_offset/$exit
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_base_plus_offset/$entry
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_base_plus_offset/sum_rename_ack
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_base_plus_offset/sum_rename_req
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_base_plus_offset/$exit
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_base_plus_offset/$entry
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_base_addr_resize/base_resize_ack
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_base_addr_resize/base_resize_ack
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_base_addr_resize/base_resize_req
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_base_addr_resize/$exit
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_base_addr_resize/$entry
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_base_addr_resize/base_resize_req
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_base_address_resized
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_root_address_calculated
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_word_address_calculated
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_base_addr_resize/$exit
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_base_address_calculated
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_base_addr_resize/$entry
      -- 
    ack_1146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_389_final_reg_ack_1, ack => testConfigure_CP_0_elements(101)); -- 
    rr_1184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(101), ack => ptr_deref_392_store_0_req_0); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	115 
    -- CP-element group 102:  members (5) 
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_Sample/word_access_start/word_0/ra
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_Sample/word_access_start/word_0/$exit
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_Sample/word_access_start/$exit
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_Sample/$exit
      -- 
    ra_1185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_392_store_0_ack_0, ack => testConfigure_CP_0_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	376 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	116 
    -- CP-element group 103:  members (5) 
      -- CP-element group 103: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_Update/word_access_complete/word_0/ca
      -- CP-element group 103: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_Update/word_access_complete/word_0/$exit
      -- CP-element group 103: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_Update/word_access_complete/$exit
      -- CP-element group 103: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_Update/$exit
      -- 
    ca_1196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_392_store_0_ack_1, ack => testConfigure_CP_0_elements(103)); -- 
    -- CP-element group 104:  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	376 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (6) 
      -- CP-element group 104: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_402_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_402_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_402_Sample/ra
      -- CP-element group 104: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_402_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_402_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_402_update_start_
      -- 
    ra_1205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_402_inst_ack_0, ack => testConfigure_CP_0_elements(104)); -- 
    cr_1209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(104), ack => RPIPE_ConvTranspose_input_pipe_402_inst_req_1); -- 
    -- CP-element group 105:  fork  transition  input  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105: 	111 
    -- CP-element group 105:  members (9) 
      -- CP-element group 105: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_418_Sample/rr
      -- CP-element group 105: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_418_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_418_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_402_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_406_Sample/rr
      -- CP-element group 105: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_406_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_406_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_402_Update/ca
      -- CP-element group 105: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_402_update_completed_
      -- 
    ca_1210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_402_inst_ack_1, ack => testConfigure_CP_0_elements(105)); -- 
    rr_1218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(105), ack => type_cast_406_inst_req_0); -- 
    rr_1282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(105), ack => RPIPE_ConvTranspose_input_pipe_418_inst_req_0); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_406_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_406_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_406_sample_completed_
      -- 
    ra_1219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_406_inst_ack_0, ack => testConfigure_CP_0_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	376 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_406_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_406_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_406_update_completed_
      -- 
    ca_1224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_406_inst_ack_1, ack => testConfigure_CP_0_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	101 
    -- CP-element group 108: 	107 
    -- CP-element group 108: 	115 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (9) 
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_Sample/word_access_start/word_0/rr
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_Sample/word_access_start/word_0/$entry
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_Sample/word_access_start/$entry
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_Sample/ptr_deref_414_Split/split_ack
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_Sample/ptr_deref_414_Split/split_req
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_Sample/ptr_deref_414_Split/$exit
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_Sample/ptr_deref_414_Split/$entry
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_Sample/$entry
      -- 
    rr_1262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(108), ack => ptr_deref_414_store_0_req_0); -- 
    testConfigure_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(101) & testConfigure_CP_0_elements(107) & testConfigure_CP_0_elements(115);
      gj_testConfigure_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (5) 
      -- CP-element group 109: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_Sample/word_access_start/word_0/ra
      -- CP-element group 109: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_Sample/word_access_start/word_0/$exit
      -- CP-element group 109: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_Sample/word_access_start/$exit
      -- CP-element group 109: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_Sample/$exit
      -- 
    ra_1263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_414_store_0_ack_0, ack => testConfigure_CP_0_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	376 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	116 
    -- CP-element group 110:  members (5) 
      -- CP-element group 110: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_Update/word_access_complete/word_0/ca
      -- CP-element group 110: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_Update/word_access_complete/word_0/$exit
      -- CP-element group 110: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_Update/word_access_complete/$exit
      -- CP-element group 110: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_Update/$exit
      -- 
    ca_1274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_414_store_0_ack_1, ack => testConfigure_CP_0_elements(110)); -- 
    -- CP-element group 111:  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	105 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (6) 
      -- CP-element group 111: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_418_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_418_Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_418_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_418_update_start_
      -- CP-element group 111: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_418_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_418_Update/cr
      -- 
    ra_1283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_418_inst_ack_0, ack => testConfigure_CP_0_elements(111)); -- 
    cr_1287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(111), ack => RPIPE_ConvTranspose_input_pipe_418_inst_req_1); -- 
    -- CP-element group 112:  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (6) 
      -- CP-element group 112: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_418_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_418_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_422_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_422_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_422_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_418_Update/ca
      -- 
    ca_1288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_418_inst_ack_1, ack => testConfigure_CP_0_elements(112)); -- 
    rr_1296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(112), ack => type_cast_422_inst_req_0); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_422_Sample/ra
      -- CP-element group 113: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_422_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_422_sample_completed_
      -- 
    ra_1297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_422_inst_ack_0, ack => testConfigure_CP_0_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	376 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_422_Update/ca
      -- CP-element group 114: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_422_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_422_update_completed_
      -- 
    ca_1302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_422_inst_ack_1, ack => testConfigure_CP_0_elements(114)); -- 
    -- CP-element group 115:  transition  delay-element  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	102 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	108 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_ptr_deref_414_delay
      -- 
    -- Element group testConfigure_CP_0_elements(115) is a control-delay.
    cp_element_115_delay: control_delay_element  generic map(name => " 115_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(102), ack => testConfigure_CP_0_elements(115), clk => clk, reset =>reset);
    -- CP-element group 116:  branch  join  transition  place  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	103 
    -- CP-element group 116: 	110 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (10) 
      -- CP-element group 116: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435__exit__
      -- CP-element group 116: 	 branch_block_stmt_34/if_stmt_436__entry__
      -- CP-element group 116: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/$exit
      -- CP-element group 116: 	 branch_block_stmt_34/R_exitcond7_437_place
      -- CP-element group 116: 	 branch_block_stmt_34/if_stmt_436_eval_test/branch_req
      -- CP-element group 116: 	 branch_block_stmt_34/if_stmt_436_eval_test/$exit
      -- CP-element group 116: 	 branch_block_stmt_34/if_stmt_436_eval_test/$entry
      -- CP-element group 116: 	 branch_block_stmt_34/if_stmt_436_dead_link/$entry
      -- CP-element group 116: 	 branch_block_stmt_34/if_stmt_436_else_link/$entry
      -- CP-element group 116: 	 branch_block_stmt_34/if_stmt_436_if_link/$entry
      -- 
    branch_req_1311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(116), ack => if_stmt_436_branch_req_0); -- 
    testConfigure_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(103) & testConfigure_CP_0_elements(110) & testConfigure_CP_0_elements(114);
      gj_testConfigure_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  fork  transition  place  input  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	377 
    -- CP-element group 117: 	378 
    -- CP-element group 117: 	380 
    -- CP-element group 117: 	381 
    -- CP-element group 117:  members (20) 
      -- CP-element group 117: 	 branch_block_stmt_34/forx_xbody69_forx_xend91
      -- CP-element group 117: 	 branch_block_stmt_34/if_stmt_436_if_link/if_choice_transition
      -- CP-element group 117: 	 branch_block_stmt_34/if_stmt_436_if_link/$exit
      -- CP-element group 117: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/$entry
      -- CP-element group 117: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_443/$entry
      -- CP-element group 117: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_443/phi_stmt_443_sources/$entry
      -- CP-element group 117: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_443/phi_stmt_443_sources/type_cast_446/$entry
      -- CP-element group 117: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_443/phi_stmt_443_sources/type_cast_446/SplitProtocol/$entry
      -- CP-element group 117: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_443/phi_stmt_443_sources/type_cast_446/SplitProtocol/Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_443/phi_stmt_443_sources/type_cast_446/SplitProtocol/Sample/rr
      -- CP-element group 117: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_443/phi_stmt_443_sources/type_cast_446/SplitProtocol/Update/$entry
      -- CP-element group 117: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_443/phi_stmt_443_sources/type_cast_446/SplitProtocol/Update/cr
      -- CP-element group 117: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_447/$entry
      -- CP-element group 117: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_447/phi_stmt_447_sources/$entry
      -- CP-element group 117: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_447/phi_stmt_447_sources/type_cast_450/$entry
      -- CP-element group 117: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_447/phi_stmt_447_sources/type_cast_450/SplitProtocol/$entry
      -- CP-element group 117: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_447/phi_stmt_447_sources/type_cast_450/SplitProtocol/Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_447/phi_stmt_447_sources/type_cast_450/SplitProtocol/Sample/rr
      -- CP-element group 117: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_447/phi_stmt_447_sources/type_cast_450/SplitProtocol/Update/$entry
      -- CP-element group 117: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_447/phi_stmt_447_sources/type_cast_450/SplitProtocol/Update/cr
      -- 
    if_choice_transition_1316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_436_branch_ack_1, ack => testConfigure_CP_0_elements(117)); -- 
    rr_3848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(117), ack => type_cast_446_inst_req_0); -- 
    cr_3853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(117), ack => type_cast_446_inst_req_1); -- 
    rr_3871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(117), ack => type_cast_450_inst_req_0); -- 
    cr_3876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(117), ack => type_cast_450_inst_req_1); -- 
    -- CP-element group 118:  fork  transition  place  input  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	366 
    -- CP-element group 118: 	367 
    -- CP-element group 118: 	369 
    -- CP-element group 118: 	370 
    -- CP-element group 118:  members (20) 
      -- CP-element group 118: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69
      -- CP-element group 118: 	 branch_block_stmt_34/if_stmt_436_else_link/else_choice_transition
      -- CP-element group 118: 	 branch_block_stmt_34/if_stmt_436_else_link/$exit
      -- CP-element group 118: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/$entry
      -- CP-element group 118: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_372/$entry
      -- CP-element group 118: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_372/phi_stmt_372_sources/$entry
      -- CP-element group 118: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_372/phi_stmt_372_sources/type_cast_378/$entry
      -- CP-element group 118: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_372/phi_stmt_372_sources/type_cast_378/SplitProtocol/$entry
      -- CP-element group 118: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_372/phi_stmt_372_sources/type_cast_378/SplitProtocol/Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_372/phi_stmt_372_sources/type_cast_378/SplitProtocol/Sample/rr
      -- CP-element group 118: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_372/phi_stmt_372_sources/type_cast_378/SplitProtocol/Update/$entry
      -- CP-element group 118: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_372/phi_stmt_372_sources/type_cast_378/SplitProtocol/Update/cr
      -- CP-element group 118: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_379/$entry
      -- CP-element group 118: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/$entry
      -- CP-element group 118: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_384/$entry
      -- CP-element group 118: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_384/SplitProtocol/$entry
      -- CP-element group 118: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_384/SplitProtocol/Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_384/SplitProtocol/Sample/rr
      -- CP-element group 118: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_384/SplitProtocol/Update/$entry
      -- CP-element group 118: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_384/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_436_branch_ack_0, ack => testConfigure_CP_0_elements(118)); -- 
    rr_3789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(118), ack => type_cast_378_inst_req_0); -- 
    cr_3794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(118), ack => type_cast_378_inst_req_1); -- 
    rr_3812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(118), ack => type_cast_384_inst_req_0); -- 
    cr_3817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(118), ack => type_cast_384_inst_req_1); -- 
    -- CP-element group 119:  join  fork  transition  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	1 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119: 	121 
    -- CP-element group 119: 	122 
    -- CP-element group 119: 	123 
    -- CP-element group 119: 	124 
    -- CP-element group 119: 	127 
    -- CP-element group 119: 	128 
    -- CP-element group 119: 	130 
    -- CP-element group 119: 	134 
    -- CP-element group 119: 	135 
    -- CP-element group 119: 	137 
    -- CP-element group 119: 	141 
    -- CP-element group 119: 	142 
    -- CP-element group 119: 	144 
    -- CP-element group 119: 	148 
    -- CP-element group 119: 	149 
    -- CP-element group 119: 	151 
    -- CP-element group 119: 	155 
    -- CP-element group 119: 	156 
    -- CP-element group 119: 	158 
    -- CP-element group 119: 	162 
    -- CP-element group 119: 	163 
    -- CP-element group 119: 	165 
    -- CP-element group 119: 	169 
    -- CP-element group 119: 	170 
    -- CP-element group 119: 	172 
    -- CP-element group 119: 	173 
    -- CP-element group 119: 	174 
    -- CP-element group 119: 	176 
    -- CP-element group 119: 	177 
    -- CP-element group 119: 	178 
    -- CP-element group 119: 	180 
    -- CP-element group 119: 	181 
    -- CP-element group 119: 	182 
    -- CP-element group 119: 	184 
    -- CP-element group 119: 	185 
    -- CP-element group 119: 	186 
    -- CP-element group 119: 	188 
    -- CP-element group 119: 	189 
    -- CP-element group 119: 	190 
    -- CP-element group 119: 	192 
    -- CP-element group 119: 	193 
    -- CP-element group 119: 	194 
    -- CP-element group 119: 	196 
    -- CP-element group 119: 	197 
    -- CP-element group 119: 	198 
    -- CP-element group 119: 	200 
    -- CP-element group 119:  members (383) 
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_root_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_base_address_resized
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_base_addr_resize/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_base_addr_resize/base_resize_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_root_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_word_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_word_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_Sample/word_access_start/word_0/rr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_word_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_Update/word_access_complete/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_Update/word_access_complete/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_Update/word_access_complete/word_0/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_base_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_base_addr_resize/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_base_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_457_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_root_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_base_address_resized
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_457_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_base_plus_offset/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_Update/word_access_complete/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_word_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_base_addr_resize/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_485_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_word_addrgen/root_register_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_731_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_457_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_base_addr_resize/base_resize_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_word_addrgen/root_register_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_base_plus_offset/sum_rename_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_base_plus_offset/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_word_addrgen/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_root_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_word_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_base_addr_resize/base_resize_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_word_addrgen/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_Update/word_access_complete/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_base_addr_resize/base_resize_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_word_addrgen/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_Update/word_access_complete/word_0/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_base_address_resized
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_457_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_base_addr_resize/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_Update/word_access_complete/word_0/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_base_addr_resize/base_resize_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_Update/word_access_complete/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_base_plus_offset/sum_rename_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_466_Sample/rr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_base_plus_offset/sum_rename_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_base_plus_offset/sum_rename_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_466_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_root_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_Update/word_access_complete/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_base_plus_offset/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_470_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_Update/word_access_complete/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_Update/word_access_complete/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_base_plus_offset/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_base_addr_resize/base_resize_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_base_plus_offset/sum_rename_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_base_addr_resize/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_base_addr_resize/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_470_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_Sample/STORE_padding_452_Split/split_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_base_plus_offset/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_Sample/STORE_padding_452_Split/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_base_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_Sample/STORE_padding_452_Split/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_457_Sample/rr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_466_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_Sample/word_access_start/word_0/rr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_base_plus_offset/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_485_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_Sample/word_access_start/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_Update/word_access_complete/word_0/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_470_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_457_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_Sample/word_access_start/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_485_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_Sample/STORE_padding_452_Split/split_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_word_addrgen/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_base_plus_offset/sum_rename_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_word_addrgen/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_word_addrgen/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_731_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_word_addrgen/root_register_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_word_addrgen/root_register_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_word_addrgen/root_register_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_word_addrgen/root_register_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_731_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_510_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_510_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_510_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_base_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_word_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_root_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_base_address_resized
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_base_addr_resize/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_base_addr_resize/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_base_addr_resize/base_resize_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_base_addr_resize/base_resize_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_base_plus_offset/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_base_plus_offset/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_base_plus_offset/sum_rename_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_base_plus_offset/sum_rename_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_word_addrgen/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_word_addrgen/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_word_addrgen/root_register_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_word_addrgen/root_register_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_Update/word_access_complete/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_Update/word_access_complete/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_Update/word_access_complete/word_0/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_534_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_534_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_534_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_base_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_word_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_root_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_base_address_resized
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_base_addr_resize/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_base_addr_resize/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_base_addr_resize/base_resize_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_base_addr_resize/base_resize_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_base_plus_offset/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_base_plus_offset/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_base_plus_offset/sum_rename_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_base_plus_offset/sum_rename_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_word_addrgen/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_word_addrgen/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_word_addrgen/root_register_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_word_addrgen/root_register_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_Sample/word_access_start/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_Update/word_access_complete/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_Update/word_access_complete/word_0/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_Update/word_access_complete/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_Update/word_access_complete/word_0/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_747_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_747_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_559_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_559_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_559_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_base_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_word_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_root_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_base_address_resized
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_base_addr_resize/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_base_addr_resize/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_base_addr_resize/base_resize_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_base_addr_resize/base_resize_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_base_plus_offset/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_base_plus_offset/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_base_plus_offset/sum_rename_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_base_plus_offset/sum_rename_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_word_addrgen/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_word_addrgen/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_word_addrgen/root_register_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_word_addrgen/root_register_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_Update/word_access_complete/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_Update/word_access_complete/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_Update/word_access_complete/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_Update/word_access_complete/word_0/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_747_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_715_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_715_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_583_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_583_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_583_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_base_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_word_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_root_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_base_address_resized
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_base_addr_resize/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_base_addr_resize/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_base_addr_resize/base_resize_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_base_addr_resize/base_resize_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_base_plus_offset/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_base_plus_offset/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_base_plus_offset/sum_rename_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_base_plus_offset/sum_rename_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_word_addrgen/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_word_addrgen/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_word_addrgen/root_register_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_word_addrgen/root_register_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_Update/word_access_complete/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_Update/word_access_complete/word_0/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_Sample/word_access_start/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_Update/word_access_complete/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_Update/word_access_complete/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_Update/word_access_complete/word_0/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_699_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_Update/word_access_complete/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_608_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_Update/word_access_complete/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_608_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_608_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_base_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_word_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_root_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_base_address_resized
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_base_addr_resize/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_base_addr_resize/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_base_addr_resize/base_resize_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_base_addr_resize/base_resize_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_base_plus_offset/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_base_plus_offset/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_base_plus_offset/sum_rename_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_base_plus_offset/sum_rename_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_word_addrgen/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_word_addrgen/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_word_addrgen/root_register_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_word_addrgen/root_register_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_Sample/word_access_start/word_0/rr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_Sample/word_access_start/word_0/rr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_699_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_Update/word_access_complete/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_Update/word_access_complete/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_Update/word_access_complete/word_0/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_Sample/word_access_start/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_715_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_Sample/word_access_start/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_base_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_word_addrgen/root_register_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_word_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_word_addrgen/root_register_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_root_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_word_addrgen/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_base_address_resized
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_base_addr_resize/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_base_addr_resize/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_base_addr_resize/base_resize_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_base_addr_resize/base_resize_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_word_addrgen/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_base_plus_offset/sum_rename_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_base_plus_offset/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_base_plus_offset/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_base_plus_offset/sum_rename_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_base_plus_offset/sum_rename_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_base_plus_offset/sum_rename_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_base_plus_offset/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_word_addrgen/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_word_addrgen/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_word_addrgen/root_register_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_word_addrgen/root_register_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_base_plus_offset/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_Sample/word_access_start/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_Sample/word_access_start/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_Sample/word_access_start/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_Sample/word_access_start/word_0/rr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_base_addr_resize/base_resize_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_Update/word_access_complete/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_Sample/word_access_start/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_Update/word_access_complete/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_Update/word_access_complete/word_0/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_base_addr_resize/base_resize_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_base_addr_resize/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_base_addr_resize/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_base_address_resized
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_641_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_root_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_641_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_641_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_word_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_base_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_base_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_word_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_root_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_base_address_resized
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_base_addr_resize/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_base_addr_resize/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_base_addr_resize/base_resize_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_base_addr_resize/base_resize_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_base_plus_offset/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_base_plus_offset/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_base_plus_offset/sum_rename_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_base_plus_offset/sum_rename_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_word_addrgen/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_word_addrgen/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_word_addrgen/root_register_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_word_addrgen/root_register_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_Sample/word_access_start/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_Sample/word_access_start/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_Sample/word_access_start/word_0/rr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_Update/word_access_complete/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_Update/word_access_complete/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_Update/word_access_complete/word_0/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_657_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_657_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_657_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_base_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_word_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_root_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_base_address_resized
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_base_addr_resize/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_base_addr_resize/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_base_addr_resize/base_resize_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_base_addr_resize/base_resize_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_base_plus_offset/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_base_plus_offset/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_base_plus_offset/sum_rename_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_base_plus_offset/sum_rename_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_word_addrgen/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_word_addrgen/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_word_addrgen/root_register_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_word_addrgen/root_register_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_Sample/word_access_start/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_Sample/word_access_start/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_Sample/word_access_start/word_0/rr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_Update/word_access_complete/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_Update/word_access_complete/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_Update/word_access_complete/word_0/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_673_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_673_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_673_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_update_start_
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_base_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_word_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_root_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_base_address_resized
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_base_addr_resize/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_base_addr_resize/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_base_addr_resize/base_resize_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_base_addr_resize/base_resize_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_base_plus_offset/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_base_plus_offset/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_base_plus_offset/sum_rename_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_base_plus_offset/sum_rename_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_word_addrgen/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_word_addrgen/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_word_addrgen/root_register_req
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_word_addrgen/root_register_ack
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_Sample/word_access_start/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_Sample/word_access_start/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_Sample/word_access_start/word_0/rr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_Update/word_access_complete/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_Update/word_access_complete/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_Update/word_access_complete/word_0/cr
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_699_update_start_
      -- 
    cr_1357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => STORE_padding_452_store_0_req_1); -- 
    rr_1346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => STORE_padding_452_store_0_req_0); -- 
    rr_1366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => type_cast_457_inst_req_0); -- 
    cr_1371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => type_cast_457_inst_req_1); -- 
    rr_1380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => RPIPE_ConvTranspose_input_pipe_466_inst_req_0); -- 
    cr_1399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => type_cast_470_inst_req_1); -- 
    cr_1432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => STORE_padding_477_store_0_req_1); -- 
    cr_1460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => type_cast_485_inst_req_1); -- 
    cr_1510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => ptr_deref_496_store_0_req_1); -- 
    cr_1538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => type_cast_510_inst_req_1); -- 
    cr_1588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => ptr_deref_526_store_0_req_1); -- 
    cr_1616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => type_cast_534_inst_req_1); -- 
    cr_1666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => ptr_deref_545_store_0_req_1); -- 
    cr_1694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => type_cast_559_inst_req_1); -- 
    cr_1744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => ptr_deref_575_store_0_req_1); -- 
    cr_1772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => type_cast_583_inst_req_1); -- 
    cr_1822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => ptr_deref_594_store_0_req_1); -- 
    cr_1850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => type_cast_608_inst_req_1); -- 
    cr_1900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => ptr_deref_624_store_0_req_1); -- 
    cr_1945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => ptr_deref_637_load_0_req_1); -- 
    rr_1934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => ptr_deref_637_load_0_req_0); -- 
    cr_1964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => type_cast_641_inst_req_1); -- 
    cr_2009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => ptr_deref_653_load_0_req_1); -- 
    rr_1998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => ptr_deref_653_load_0_req_0); -- 
    cr_2028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => type_cast_657_inst_req_1); -- 
    cr_2073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => ptr_deref_669_load_0_req_1); -- 
    rr_2062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => ptr_deref_669_load_0_req_0); -- 
    cr_2092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => type_cast_673_inst_req_1); -- 
    cr_2137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => ptr_deref_695_load_0_req_1); -- 
    rr_2126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => ptr_deref_695_load_0_req_0); -- 
    cr_2156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => type_cast_699_inst_req_1); -- 
    cr_2201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => ptr_deref_711_load_0_req_1); -- 
    rr_2190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => ptr_deref_711_load_0_req_0); -- 
    cr_2220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => type_cast_715_inst_req_1); -- 
    cr_2265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => ptr_deref_727_load_0_req_1); -- 
    rr_2254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => ptr_deref_727_load_0_req_0); -- 
    cr_2284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => type_cast_731_inst_req_1); -- 
    cr_2329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => ptr_deref_743_load_0_req_1); -- 
    rr_2318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => ptr_deref_743_load_0_req_0); -- 
    cr_2348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => type_cast_747_inst_req_1); -- 
    testConfigure_CP_0_elements(119) <= testConfigure_CP_0_elements(1);
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	206 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_Sample/word_access_start/$exit
      -- CP-element group 120: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_Sample/word_access_start/word_0/ra
      -- CP-element group 120: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_Sample/word_access_start/word_0/$exit
      -- CP-element group 120: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_Sample/$exit
      -- 
    ra_1347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_padding_452_store_0_ack_0, ack => testConfigure_CP_0_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	207 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_Update/word_access_complete/word_0/ca
      -- CP-element group 121: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_Update/word_access_complete/word_0/$exit
      -- CP-element group 121: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_Update/word_access_complete/$exit
      -- CP-element group 121: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_Update/$exit
      -- 
    ca_1358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_padding_452_store_0_ack_1, ack => testConfigure_CP_0_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	119 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_457_sample_completed_
      -- CP-element group 122: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_457_Sample/$exit
      -- CP-element group 122: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_457_Sample/ra
      -- 
    ra_1367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_457_inst_ack_0, ack => testConfigure_CP_0_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	119 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	128 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_457_Update/ca
      -- CP-element group 123: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_457_Update/$exit
      -- CP-element group 123: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_457_update_completed_
      -- 
    ca_1372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_457_inst_ack_1, ack => testConfigure_CP_0_elements(123)); -- 
    -- CP-element group 124:  transition  input  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	119 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (6) 
      -- CP-element group 124: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_466_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_466_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_466_Sample/ra
      -- CP-element group 124: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_466_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_466_update_start_
      -- CP-element group 124: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_466_sample_completed_
      -- 
    ra_1381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_466_inst_ack_0, ack => testConfigure_CP_0_elements(124)); -- 
    cr_1385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(124), ack => RPIPE_ConvTranspose_input_pipe_466_inst_req_1); -- 
    -- CP-element group 125:  fork  transition  input  output  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125: 	131 
    -- CP-element group 125:  members (9) 
      -- CP-element group 125: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_470_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_481_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_466_Update/ca
      -- CP-element group 125: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_466_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_466_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_481_Sample/rr
      -- CP-element group 125: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_470_Sample/rr
      -- CP-element group 125: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_470_Sample/$entry
      -- CP-element group 125: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_481_Sample/$entry
      -- 
    ca_1386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_466_inst_ack_1, ack => testConfigure_CP_0_elements(125)); -- 
    rr_1394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(125), ack => type_cast_470_inst_req_0); -- 
    rr_1441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(125), ack => RPIPE_ConvTranspose_input_pipe_481_inst_req_0); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_470_Sample/ra
      -- CP-element group 126: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_470_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_470_sample_completed_
      -- 
    ra_1395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_470_inst_ack_0, ack => testConfigure_CP_0_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	119 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_470_Update/ca
      -- CP-element group 127: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_470_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_470_update_completed_
      -- 
    ca_1400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_470_inst_ack_1, ack => testConfigure_CP_0_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	119 
    -- CP-element group 128: 	123 
    -- CP-element group 128: 	127 
    -- CP-element group 128: 	206 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (9) 
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_Sample/word_access_start/$entry
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_Sample/STORE_padding_477_Split/split_ack
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_Sample/STORE_padding_477_Split/split_req
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_Sample/STORE_padding_477_Split/$exit
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_Sample/STORE_padding_477_Split/$entry
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_Sample/word_access_start/word_0/rr
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_Sample/word_access_start/word_0/$entry
      -- 
    rr_1421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(128), ack => STORE_padding_477_store_0_req_0); -- 
    testConfigure_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(119) & testConfigure_CP_0_elements(123) & testConfigure_CP_0_elements(127) & testConfigure_CP_0_elements(206);
      gj_testConfigure_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (5) 
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_Sample/word_access_start/$exit
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_Sample/word_access_start/word_0/ra
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_Sample/word_access_start/word_0/$exit
      -- 
    ra_1422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_padding_477_store_0_ack_0, ack => testConfigure_CP_0_elements(129)); -- 
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	119 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	207 
    -- CP-element group 130:  members (5) 
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_Update/word_access_complete/word_0/ca
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_Update/word_access_complete/word_0/$exit
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_Update/word_access_complete/$exit
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_477_Update/$exit
      -- 
    ca_1433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_padding_477_store_0_ack_1, ack => testConfigure_CP_0_elements(130)); -- 
    -- CP-element group 131:  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	125 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (6) 
      -- CP-element group 131: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_481_update_start_
      -- CP-element group 131: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_481_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_481_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_481_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_481_Sample/ra
      -- CP-element group 131: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_481_Sample/$exit
      -- 
    ra_1442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_481_inst_ack_0, ack => testConfigure_CP_0_elements(131)); -- 
    cr_1446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(131), ack => RPIPE_ConvTranspose_input_pipe_481_inst_req_1); -- 
    -- CP-element group 132:  fork  transition  input  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132: 	138 
    -- CP-element group 132:  members (9) 
      -- CP-element group 132: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_506_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_506_Sample/rr
      -- CP-element group 132: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_506_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_481_Update/ca
      -- CP-element group 132: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_481_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_481_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_485_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_485_Sample/rr
      -- CP-element group 132: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_485_Sample/$entry
      -- 
    ca_1447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_481_inst_ack_1, ack => testConfigure_CP_0_elements(132)); -- 
    rr_1455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(132), ack => type_cast_485_inst_req_0); -- 
    rr_1519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(132), ack => RPIPE_ConvTranspose_input_pipe_506_inst_req_0); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_485_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_485_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_485_Sample/$exit
      -- 
    ra_1456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_485_inst_ack_0, ack => testConfigure_CP_0_elements(133)); -- 
    -- CP-element group 134:  fork  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	119 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	142 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_485_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_485_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_485_Update/ca
      -- 
    ca_1461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_485_inst_ack_1, ack => testConfigure_CP_0_elements(134)); -- 
    -- CP-element group 135:  join  transition  output  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	119 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (9) 
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_Sample/ptr_deref_496_Split/split_ack
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_Sample/word_access_start/$entry
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_Sample/word_access_start/word_0/$entry
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_Sample/word_access_start/word_0/rr
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_Sample/ptr_deref_496_Split/split_req
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_Sample/ptr_deref_496_Split/$entry
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_Sample/ptr_deref_496_Split/$exit
      -- 
    rr_1499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(135), ack => ptr_deref_496_store_0_req_0); -- 
    testConfigure_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(119) & testConfigure_CP_0_elements(134);
      gj_testConfigure_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	201 
    -- CP-element group 136:  members (5) 
      -- CP-element group 136: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_Sample/word_access_start/word_0/ra
      -- CP-element group 136: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_Sample/word_access_start/word_0/$exit
      -- CP-element group 136: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_Sample/word_access_start/$exit
      -- CP-element group 136: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_Sample/$exit
      -- 
    ra_1500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_496_store_0_ack_0, ack => testConfigure_CP_0_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	119 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	207 
    -- CP-element group 137:  members (5) 
      -- CP-element group 137: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_Update/word_access_complete/word_0/ca
      -- CP-element group 137: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_Update/word_access_complete/word_0/$exit
      -- CP-element group 137: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_Update/word_access_complete/$exit
      -- CP-element group 137: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_Update/$exit
      -- 
    ca_1511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_496_store_0_ack_1, ack => testConfigure_CP_0_elements(137)); -- 
    -- CP-element group 138:  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	132 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138:  members (6) 
      -- CP-element group 138: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_506_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_506_Sample/ra
      -- CP-element group 138: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_506_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_506_sample_completed_
      -- CP-element group 138: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_506_update_start_
      -- CP-element group 138: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_506_Update/cr
      -- 
    ra_1520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_506_inst_ack_0, ack => testConfigure_CP_0_elements(138)); -- 
    cr_1524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(138), ack => RPIPE_ConvTranspose_input_pipe_506_inst_req_1); -- 
    -- CP-element group 139:  fork  transition  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	140 
    -- CP-element group 139: 	145 
    -- CP-element group 139:  members (9) 
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_506_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_506_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_506_Update/ca
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_510_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_510_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_510_Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_530_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_530_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_530_Sample/rr
      -- 
    ca_1525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_506_inst_ack_1, ack => testConfigure_CP_0_elements(139)); -- 
    rr_1533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(139), ack => type_cast_510_inst_req_0); -- 
    rr_1597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(139), ack => RPIPE_ConvTranspose_input_pipe_530_inst_req_0); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	139 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_510_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_510_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_510_Sample/ra
      -- 
    ra_1534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_510_inst_ack_0, ack => testConfigure_CP_0_elements(140)); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	119 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_510_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_510_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_510_Update/ca
      -- 
    ca_1539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_510_inst_ack_1, ack => testConfigure_CP_0_elements(141)); -- 
    -- CP-element group 142:  join  transition  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	119 
    -- CP-element group 142: 	134 
    -- CP-element group 142: 	141 
    -- CP-element group 142: 	201 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142:  members (9) 
      -- CP-element group 142: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_Sample/ptr_deref_526_Split/$entry
      -- CP-element group 142: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_Sample/ptr_deref_526_Split/$exit
      -- CP-element group 142: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_Sample/ptr_deref_526_Split/split_req
      -- CP-element group 142: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_Sample/ptr_deref_526_Split/split_ack
      -- CP-element group 142: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_Sample/word_access_start/$entry
      -- CP-element group 142: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_Sample/word_access_start/word_0/$entry
      -- CP-element group 142: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_Sample/word_access_start/word_0/rr
      -- 
    rr_1577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(142), ack => ptr_deref_526_store_0_req_0); -- 
    testConfigure_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(119) & testConfigure_CP_0_elements(134) & testConfigure_CP_0_elements(141) & testConfigure_CP_0_elements(201);
      gj_testConfigure_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	202 
    -- CP-element group 143:  members (5) 
      -- CP-element group 143: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_Sample/word_access_start/$exit
      -- CP-element group 143: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_Sample/word_access_start/word_0/$exit
      -- CP-element group 143: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_Sample/word_access_start/word_0/ra
      -- 
    ra_1578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_526_store_0_ack_0, ack => testConfigure_CP_0_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	119 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	207 
    -- CP-element group 144:  members (5) 
      -- CP-element group 144: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_Update/word_access_complete/$exit
      -- CP-element group 144: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_Update/word_access_complete/word_0/$exit
      -- CP-element group 144: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_Update/word_access_complete/word_0/ca
      -- 
    ca_1589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_526_store_0_ack_1, ack => testConfigure_CP_0_elements(144)); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	139 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_530_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_530_update_start_
      -- CP-element group 145: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_530_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_530_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_530_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_530_Update/cr
      -- 
    ra_1598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_530_inst_ack_0, ack => testConfigure_CP_0_elements(145)); -- 
    cr_1602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(145), ack => RPIPE_ConvTranspose_input_pipe_530_inst_req_1); -- 
    -- CP-element group 146:  fork  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	152 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_530_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_530_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_530_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_534_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_534_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_534_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_555_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_555_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_555_Sample/rr
      -- 
    ca_1603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_530_inst_ack_1, ack => testConfigure_CP_0_elements(146)); -- 
    rr_1611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(146), ack => type_cast_534_inst_req_0); -- 
    rr_1675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(146), ack => RPIPE_ConvTranspose_input_pipe_555_inst_req_0); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_534_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_534_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_534_Sample/ra
      -- 
    ra_1612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_534_inst_ack_0, ack => testConfigure_CP_0_elements(147)); -- 
    -- CP-element group 148:  fork  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	119 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: 	156 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_534_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_534_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_534_Update/ca
      -- 
    ca_1617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_534_inst_ack_1, ack => testConfigure_CP_0_elements(148)); -- 
    -- CP-element group 149:  join  transition  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	119 
    -- CP-element group 149: 	148 
    -- CP-element group 149: 	202 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (9) 
      -- CP-element group 149: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_sample_start_
      -- CP-element group 149: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_Sample/ptr_deref_545_Split/$entry
      -- CP-element group 149: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_Sample/ptr_deref_545_Split/$exit
      -- CP-element group 149: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_Sample/ptr_deref_545_Split/split_req
      -- CP-element group 149: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_Sample/ptr_deref_545_Split/split_ack
      -- CP-element group 149: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_Sample/word_access_start/$entry
      -- CP-element group 149: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_Sample/word_access_start/word_0/$entry
      -- CP-element group 149: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_Sample/word_access_start/word_0/rr
      -- 
    rr_1655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(149), ack => ptr_deref_545_store_0_req_0); -- 
    testConfigure_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(119) & testConfigure_CP_0_elements(148) & testConfigure_CP_0_elements(202);
      gj_testConfigure_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	203 
    -- CP-element group 150:  members (5) 
      -- CP-element group 150: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_sample_completed_
      -- CP-element group 150: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_Sample/$exit
      -- CP-element group 150: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_Sample/word_access_start/$exit
      -- CP-element group 150: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_Sample/word_access_start/word_0/$exit
      -- CP-element group 150: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_Sample/word_access_start/word_0/ra
      -- 
    ra_1656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_545_store_0_ack_0, ack => testConfigure_CP_0_elements(150)); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	119 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	207 
    -- CP-element group 151:  members (5) 
      -- CP-element group 151: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_update_completed_
      -- CP-element group 151: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_Update/$exit
      -- CP-element group 151: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_Update/word_access_complete/$exit
      -- CP-element group 151: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_Update/word_access_complete/word_0/$exit
      -- CP-element group 151: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_Update/word_access_complete/word_0/ca
      -- 
    ca_1667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_545_store_0_ack_1, ack => testConfigure_CP_0_elements(151)); -- 
    -- CP-element group 152:  transition  input  output  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	146 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152:  members (6) 
      -- CP-element group 152: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_555_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_555_update_start_
      -- CP-element group 152: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_555_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_555_Sample/ra
      -- CP-element group 152: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_555_Update/$entry
      -- CP-element group 152: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_555_Update/cr
      -- 
    ra_1676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_555_inst_ack_0, ack => testConfigure_CP_0_elements(152)); -- 
    cr_1680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(152), ack => RPIPE_ConvTranspose_input_pipe_555_inst_req_1); -- 
    -- CP-element group 153:  fork  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	152 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153: 	159 
    -- CP-element group 153:  members (9) 
      -- CP-element group 153: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_555_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_555_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_555_Update/ca
      -- CP-element group 153: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_559_sample_start_
      -- CP-element group 153: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_559_Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_559_Sample/rr
      -- CP-element group 153: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_579_sample_start_
      -- CP-element group 153: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_579_Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_579_Sample/rr
      -- 
    ca_1681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_555_inst_ack_1, ack => testConfigure_CP_0_elements(153)); -- 
    rr_1689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(153), ack => type_cast_559_inst_req_0); -- 
    rr_1753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(153), ack => RPIPE_ConvTranspose_input_pipe_579_inst_req_0); -- 
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_559_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_559_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_559_Sample/ra
      -- 
    ra_1690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_559_inst_ack_0, ack => testConfigure_CP_0_elements(154)); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	119 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_559_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_559_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_559_Update/ca
      -- 
    ca_1695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_559_inst_ack_1, ack => testConfigure_CP_0_elements(155)); -- 
    -- CP-element group 156:  join  transition  output  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	119 
    -- CP-element group 156: 	148 
    -- CP-element group 156: 	155 
    -- CP-element group 156: 	203 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	157 
    -- CP-element group 156:  members (9) 
      -- CP-element group 156: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_Sample/ptr_deref_575_Split/$entry
      -- CP-element group 156: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_Sample/ptr_deref_575_Split/$exit
      -- CP-element group 156: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_Sample/ptr_deref_575_Split/split_req
      -- CP-element group 156: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_Sample/ptr_deref_575_Split/split_ack
      -- CP-element group 156: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_Sample/word_access_start/$entry
      -- CP-element group 156: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_Sample/word_access_start/word_0/$entry
      -- CP-element group 156: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_Sample/word_access_start/word_0/rr
      -- 
    rr_1733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(156), ack => ptr_deref_575_store_0_req_0); -- 
    testConfigure_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(119) & testConfigure_CP_0_elements(148) & testConfigure_CP_0_elements(155) & testConfigure_CP_0_elements(203);
      gj_testConfigure_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	156 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	204 
    -- CP-element group 157:  members (5) 
      -- CP-element group 157: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_Sample/word_access_start/$exit
      -- CP-element group 157: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_Sample/word_access_start/word_0/$exit
      -- CP-element group 157: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_Sample/word_access_start/word_0/ra
      -- 
    ra_1734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_575_store_0_ack_0, ack => testConfigure_CP_0_elements(157)); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	119 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	207 
    -- CP-element group 158:  members (5) 
      -- CP-element group 158: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_Update/word_access_complete/$exit
      -- CP-element group 158: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_Update/word_access_complete/word_0/$exit
      -- CP-element group 158: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_Update/word_access_complete/word_0/ca
      -- 
    ca_1745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_575_store_0_ack_1, ack => testConfigure_CP_0_elements(158)); -- 
    -- CP-element group 159:  transition  input  output  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	153 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159:  members (6) 
      -- CP-element group 159: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_579_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_579_update_start_
      -- CP-element group 159: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_579_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_579_Sample/ra
      -- CP-element group 159: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_579_Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_579_Update/cr
      -- 
    ra_1754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_579_inst_ack_0, ack => testConfigure_CP_0_elements(159)); -- 
    cr_1758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(159), ack => RPIPE_ConvTranspose_input_pipe_579_inst_req_1); -- 
    -- CP-element group 160:  fork  transition  input  output  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	159 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160: 	166 
    -- CP-element group 160:  members (9) 
      -- CP-element group 160: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_579_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_579_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_579_Update/ca
      -- CP-element group 160: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_583_sample_start_
      -- CP-element group 160: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_583_Sample/$entry
      -- CP-element group 160: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_583_Sample/rr
      -- CP-element group 160: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_604_sample_start_
      -- CP-element group 160: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_604_Sample/$entry
      -- CP-element group 160: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_604_Sample/rr
      -- 
    ca_1759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_579_inst_ack_1, ack => testConfigure_CP_0_elements(160)); -- 
    rr_1767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(160), ack => type_cast_583_inst_req_0); -- 
    rr_1831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(160), ack => RPIPE_ConvTranspose_input_pipe_604_inst_req_0); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_583_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_583_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_583_Sample/ra
      -- 
    ra_1768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_583_inst_ack_0, ack => testConfigure_CP_0_elements(161)); -- 
    -- CP-element group 162:  fork  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	119 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162: 	170 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_583_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_583_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_583_Update/ca
      -- 
    ca_1773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_583_inst_ack_1, ack => testConfigure_CP_0_elements(162)); -- 
    -- CP-element group 163:  join  transition  output  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	119 
    -- CP-element group 163: 	162 
    -- CP-element group 163: 	204 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (9) 
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_Sample/ptr_deref_594_Split/$entry
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_Sample/ptr_deref_594_Split/$exit
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_Sample/ptr_deref_594_Split/split_req
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_Sample/ptr_deref_594_Split/split_ack
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_Sample/word_access_start/$entry
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_Sample/word_access_start/word_0/$entry
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_Sample/word_access_start/word_0/rr
      -- 
    rr_1811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(163), ack => ptr_deref_594_store_0_req_0); -- 
    testConfigure_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(119) & testConfigure_CP_0_elements(162) & testConfigure_CP_0_elements(204);
      gj_testConfigure_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	205 
    -- CP-element group 164:  members (5) 
      -- CP-element group 164: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_sample_completed_
      -- CP-element group 164: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_Sample/word_access_start/$exit
      -- CP-element group 164: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_Sample/word_access_start/word_0/$exit
      -- CP-element group 164: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_Sample/word_access_start/word_0/ra
      -- 
    ra_1812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_594_store_0_ack_0, ack => testConfigure_CP_0_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	119 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	207 
    -- CP-element group 165:  members (5) 
      -- CP-element group 165: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_Update/word_access_complete/$exit
      -- CP-element group 165: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_Update/word_access_complete/word_0/$exit
      -- CP-element group 165: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_Update/word_access_complete/word_0/ca
      -- 
    ca_1823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_594_store_0_ack_1, ack => testConfigure_CP_0_elements(165)); -- 
    -- CP-element group 166:  transition  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	160 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166:  members (6) 
      -- CP-element group 166: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_604_sample_completed_
      -- CP-element group 166: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_604_update_start_
      -- CP-element group 166: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_604_Sample/$exit
      -- CP-element group 166: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_604_Sample/ra
      -- CP-element group 166: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_604_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_604_Update/cr
      -- 
    ra_1832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_604_inst_ack_0, ack => testConfigure_CP_0_elements(166)); -- 
    cr_1836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(166), ack => RPIPE_ConvTranspose_input_pipe_604_inst_req_1); -- 
    -- CP-element group 167:  transition  input  output  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	168 
    -- CP-element group 167:  members (6) 
      -- CP-element group 167: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_604_update_completed_
      -- CP-element group 167: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_604_Update/$exit
      -- CP-element group 167: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/RPIPE_ConvTranspose_input_pipe_604_Update/ca
      -- CP-element group 167: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_608_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_608_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_608_Sample/rr
      -- 
    ca_1837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_604_inst_ack_1, ack => testConfigure_CP_0_elements(167)); -- 
    rr_1845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(167), ack => type_cast_608_inst_req_0); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	167 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_608_sample_completed_
      -- CP-element group 168: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_608_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_608_Sample/ra
      -- 
    ra_1846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_608_inst_ack_0, ack => testConfigure_CP_0_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	119 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_608_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_608_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_608_Update/ca
      -- 
    ca_1851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_608_inst_ack_1, ack => testConfigure_CP_0_elements(169)); -- 
    -- CP-element group 170:  join  transition  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	119 
    -- CP-element group 170: 	162 
    -- CP-element group 170: 	169 
    -- CP-element group 170: 	205 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (9) 
      -- CP-element group 170: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_Sample/$entry
      -- CP-element group 170: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_Sample/ptr_deref_624_Split/$entry
      -- CP-element group 170: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_Sample/ptr_deref_624_Split/$exit
      -- CP-element group 170: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_Sample/ptr_deref_624_Split/split_req
      -- CP-element group 170: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_Sample/ptr_deref_624_Split/split_ack
      -- CP-element group 170: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_Sample/word_access_start/$entry
      -- CP-element group 170: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_Sample/word_access_start/word_0/$entry
      -- CP-element group 170: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_Sample/word_access_start/word_0/rr
      -- 
    rr_1889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(170), ack => ptr_deref_624_store_0_req_0); -- 
    testConfigure_cp_element_group_170: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_170"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(119) & testConfigure_CP_0_elements(162) & testConfigure_CP_0_elements(169) & testConfigure_CP_0_elements(205);
      gj_testConfigure_cp_element_group_170 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(170), clk => clk, reset => reset); --
    end block;
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (5) 
      -- CP-element group 171: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_Sample/word_access_start/$exit
      -- CP-element group 171: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_Sample/word_access_start/word_0/$exit
      -- CP-element group 171: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_Sample/word_access_start/word_0/ra
      -- 
    ra_1890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_624_store_0_ack_0, ack => testConfigure_CP_0_elements(171)); -- 
    -- CP-element group 172:  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	119 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	207 
    -- CP-element group 172:  members (5) 
      -- CP-element group 172: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_Update/word_access_complete/$exit
      -- CP-element group 172: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_Update/word_access_complete/word_0/$exit
      -- CP-element group 172: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_624_Update/word_access_complete/word_0/ca
      -- 
    ca_1901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_624_store_0_ack_1, ack => testConfigure_CP_0_elements(172)); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	119 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (5) 
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_Sample/word_access_start/$exit
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_Sample/word_access_start/word_0/$exit
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_Sample/word_access_start/word_0/ra
      -- 
    ra_1935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_637_load_0_ack_0, ack => testConfigure_CP_0_elements(173)); -- 
    -- CP-element group 174:  transition  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	119 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174:  members (12) 
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_Update/word_access_complete/$exit
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_Update/word_access_complete/word_0/$exit
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_Update/word_access_complete/word_0/ca
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_Update/ptr_deref_637_Merge/$entry
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_Update/ptr_deref_637_Merge/$exit
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_Update/ptr_deref_637_Merge/merge_req
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_637_Update/ptr_deref_637_Merge/merge_ack
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_641_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_641_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_641_Sample/rr
      -- 
    ca_1946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_637_load_0_ack_1, ack => testConfigure_CP_0_elements(174)); -- 
    rr_1959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(174), ack => type_cast_641_inst_req_0); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_641_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_641_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_641_Sample/ra
      -- 
    ra_1960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_641_inst_ack_0, ack => testConfigure_CP_0_elements(175)); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	119 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	207 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_641_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_641_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_641_Update/ca
      -- 
    ca_1965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_641_inst_ack_1, ack => testConfigure_CP_0_elements(176)); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	119 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (5) 
      -- CP-element group 177: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_Sample/word_access_start/$exit
      -- CP-element group 177: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_Sample/word_access_start/word_0/$exit
      -- CP-element group 177: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_Sample/word_access_start/word_0/ra
      -- 
    ra_1999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_653_load_0_ack_0, ack => testConfigure_CP_0_elements(177)); -- 
    -- CP-element group 178:  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	119 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (12) 
      -- CP-element group 178: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_Update/word_access_complete/$exit
      -- CP-element group 178: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_Update/word_access_complete/word_0/$exit
      -- CP-element group 178: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_Update/word_access_complete/word_0/ca
      -- CP-element group 178: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_Update/ptr_deref_653_Merge/$entry
      -- CP-element group 178: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_Update/ptr_deref_653_Merge/$exit
      -- CP-element group 178: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_Update/ptr_deref_653_Merge/merge_req
      -- CP-element group 178: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_653_Update/ptr_deref_653_Merge/merge_ack
      -- CP-element group 178: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_657_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_657_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_657_Sample/rr
      -- 
    ca_2010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_653_load_0_ack_1, ack => testConfigure_CP_0_elements(178)); -- 
    rr_2023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(178), ack => type_cast_657_inst_req_0); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_657_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_657_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_657_Sample/ra
      -- 
    ra_2024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_657_inst_ack_0, ack => testConfigure_CP_0_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	119 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	207 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_657_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_657_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_657_Update/ca
      -- 
    ca_2029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_657_inst_ack_1, ack => testConfigure_CP_0_elements(180)); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	119 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (5) 
      -- CP-element group 181: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_Sample/word_access_start/$exit
      -- CP-element group 181: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_Sample/word_access_start/word_0/$exit
      -- CP-element group 181: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_Sample/word_access_start/word_0/ra
      -- 
    ra_2063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_669_load_0_ack_0, ack => testConfigure_CP_0_elements(181)); -- 
    -- CP-element group 182:  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	119 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182:  members (12) 
      -- CP-element group 182: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_Update/word_access_complete/$exit
      -- CP-element group 182: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_Update/word_access_complete/word_0/$exit
      -- CP-element group 182: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_Update/word_access_complete/word_0/ca
      -- CP-element group 182: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_Update/ptr_deref_669_Merge/$entry
      -- CP-element group 182: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_Update/ptr_deref_669_Merge/$exit
      -- CP-element group 182: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_Update/ptr_deref_669_Merge/merge_req
      -- CP-element group 182: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_669_Update/ptr_deref_669_Merge/merge_ack
      -- CP-element group 182: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_673_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_673_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_673_Sample/rr
      -- 
    ca_2074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_669_load_0_ack_1, ack => testConfigure_CP_0_elements(182)); -- 
    rr_2087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(182), ack => type_cast_673_inst_req_0); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_673_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_673_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_673_Sample/ra
      -- 
    ra_2088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_673_inst_ack_0, ack => testConfigure_CP_0_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	119 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	207 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_673_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_673_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_673_Update/ca
      -- 
    ca_2093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_673_inst_ack_1, ack => testConfigure_CP_0_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	119 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (5) 
      -- CP-element group 185: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_Sample/word_access_start/$exit
      -- CP-element group 185: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_Sample/word_access_start/word_0/$exit
      -- CP-element group 185: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_Sample/word_access_start/word_0/ra
      -- 
    ra_2127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_695_load_0_ack_0, ack => testConfigure_CP_0_elements(185)); -- 
    -- CP-element group 186:  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	119 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (12) 
      -- CP-element group 186: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_699_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_699_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_Update/word_access_complete/$exit
      -- CP-element group 186: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_Update/word_access_complete/word_0/$exit
      -- CP-element group 186: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_Update/word_access_complete/word_0/ca
      -- CP-element group 186: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_Update/ptr_deref_695_Merge/$entry
      -- CP-element group 186: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_Update/ptr_deref_695_Merge/$exit
      -- CP-element group 186: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_Update/ptr_deref_695_Merge/merge_req
      -- CP-element group 186: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_695_Update/ptr_deref_695_Merge/merge_ack
      -- CP-element group 186: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_699_sample_start_
      -- 
    ca_2138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_695_load_0_ack_1, ack => testConfigure_CP_0_elements(186)); -- 
    rr_2151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(186), ack => type_cast_699_inst_req_0); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_699_Sample/ra
      -- CP-element group 187: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_699_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_699_sample_completed_
      -- 
    ra_2152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_699_inst_ack_0, ack => testConfigure_CP_0_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	119 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	207 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_699_Update/ca
      -- CP-element group 188: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_699_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_699_update_completed_
      -- 
    ca_2157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_699_inst_ack_1, ack => testConfigure_CP_0_elements(188)); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	119 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (5) 
      -- CP-element group 189: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_Sample/word_access_start/word_0/ra
      -- CP-element group 189: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_Sample/word_access_start/word_0/$exit
      -- CP-element group 189: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_Sample/word_access_start/$exit
      -- 
    ra_2191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_711_load_0_ack_0, ack => testConfigure_CP_0_elements(189)); -- 
    -- CP-element group 190:  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	119 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190:  members (12) 
      -- CP-element group 190: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_Update/word_access_complete/$exit
      -- CP-element group 190: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_Update/word_access_complete/word_0/$exit
      -- CP-element group 190: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_Update/word_access_complete/word_0/ca
      -- CP-element group 190: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_715_Sample/rr
      -- CP-element group 190: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_715_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_715_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_Update/ptr_deref_711_Merge/merge_ack
      -- CP-element group 190: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_Update/ptr_deref_711_Merge/merge_req
      -- CP-element group 190: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_Update/ptr_deref_711_Merge/$exit
      -- CP-element group 190: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_711_Update/ptr_deref_711_Merge/$entry
      -- 
    ca_2202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_711_load_0_ack_1, ack => testConfigure_CP_0_elements(190)); -- 
    rr_2215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(190), ack => type_cast_715_inst_req_0); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_715_Sample/ra
      -- CP-element group 191: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_715_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_715_sample_completed_
      -- 
    ra_2216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_715_inst_ack_0, ack => testConfigure_CP_0_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	119 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	207 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_715_Update/ca
      -- CP-element group 192: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_715_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_715_update_completed_
      -- 
    ca_2221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_715_inst_ack_1, ack => testConfigure_CP_0_elements(192)); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	119 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (5) 
      -- CP-element group 193: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_Sample/word_access_start/word_0/ra
      -- CP-element group 193: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_Sample/word_access_start/word_0/$exit
      -- CP-element group 193: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_Sample/word_access_start/$exit
      -- 
    ra_2255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_727_load_0_ack_0, ack => testConfigure_CP_0_elements(193)); -- 
    -- CP-element group 194:  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	119 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (12) 
      -- CP-element group 194: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_731_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_731_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_731_Sample/rr
      -- CP-element group 194: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_Update/ptr_deref_727_Merge/merge_ack
      -- CP-element group 194: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_Update/ptr_deref_727_Merge/merge_req
      -- CP-element group 194: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_Update/ptr_deref_727_Merge/$exit
      -- CP-element group 194: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_Update/ptr_deref_727_Merge/$entry
      -- CP-element group 194: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_Update/word_access_complete/word_0/ca
      -- CP-element group 194: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_Update/word_access_complete/word_0/$exit
      -- CP-element group 194: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_Update/word_access_complete/$exit
      -- CP-element group 194: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_727_Update/$exit
      -- 
    ca_2266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_727_load_0_ack_1, ack => testConfigure_CP_0_elements(194)); -- 
    rr_2279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(194), ack => type_cast_731_inst_req_0); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_731_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_731_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_731_Sample/ra
      -- 
    ra_2280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_731_inst_ack_0, ack => testConfigure_CP_0_elements(195)); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	119 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	207 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_731_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_731_Update/ca
      -- CP-element group 196: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_731_Update/$exit
      -- 
    ca_2285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_731_inst_ack_1, ack => testConfigure_CP_0_elements(196)); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	119 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (5) 
      -- CP-element group 197: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_Sample/word_access_start/word_0/ra
      -- CP-element group 197: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_Sample/word_access_start/word_0/$exit
      -- CP-element group 197: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_Sample/word_access_start/$exit
      -- CP-element group 197: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_sample_completed_
      -- 
    ra_2319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_743_load_0_ack_0, ack => testConfigure_CP_0_elements(197)); -- 
    -- CP-element group 198:  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	119 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198:  members (12) 
      -- CP-element group 198: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_747_Sample/rr
      -- CP-element group 198: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_747_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_747_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_Update/ptr_deref_743_Merge/merge_ack
      -- CP-element group 198: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_Update/ptr_deref_743_Merge/merge_req
      -- CP-element group 198: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_Update/ptr_deref_743_Merge/$exit
      -- CP-element group 198: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_Update/ptr_deref_743_Merge/$entry
      -- CP-element group 198: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_Update/word_access_complete/word_0/ca
      -- CP-element group 198: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_Update/word_access_complete/word_0/$exit
      -- CP-element group 198: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_Update/word_access_complete/$exit
      -- CP-element group 198: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_743_update_completed_
      -- 
    ca_2330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_743_load_0_ack_1, ack => testConfigure_CP_0_elements(198)); -- 
    rr_2343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(198), ack => type_cast_747_inst_req_0); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_747_Sample/ra
      -- CP-element group 199: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_747_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_747_sample_completed_
      -- 
    ra_2344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_747_inst_ack_0, ack => testConfigure_CP_0_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	119 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	207 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_747_Update/ca
      -- CP-element group 200: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_747_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/type_cast_747_update_completed_
      -- 
    ca_2349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_747_inst_ack_1, ack => testConfigure_CP_0_elements(200)); -- 
    -- CP-element group 201:  transition  delay-element  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	136 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	142 
    -- CP-element group 201:  members (1) 
      -- CP-element group 201: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_496_ptr_deref_526_delay
      -- 
    -- Element group testConfigure_CP_0_elements(201) is a control-delay.
    cp_element_201_delay: control_delay_element  generic map(name => " 201_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(136), ack => testConfigure_CP_0_elements(201), clk => clk, reset =>reset);
    -- CP-element group 202:  transition  delay-element  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	143 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	149 
    -- CP-element group 202:  members (1) 
      -- CP-element group 202: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_526_ptr_deref_545_delay
      -- 
    -- Element group testConfigure_CP_0_elements(202) is a control-delay.
    cp_element_202_delay: control_delay_element  generic map(name => " 202_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(143), ack => testConfigure_CP_0_elements(202), clk => clk, reset =>reset);
    -- CP-element group 203:  transition  delay-element  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	150 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	156 
    -- CP-element group 203:  members (1) 
      -- CP-element group 203: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_545_ptr_deref_575_delay
      -- 
    -- Element group testConfigure_CP_0_elements(203) is a control-delay.
    cp_element_203_delay: control_delay_element  generic map(name => " 203_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(150), ack => testConfigure_CP_0_elements(203), clk => clk, reset =>reset);
    -- CP-element group 204:  transition  delay-element  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	157 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	163 
    -- CP-element group 204:  members (1) 
      -- CP-element group 204: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_575_ptr_deref_594_delay
      -- 
    -- Element group testConfigure_CP_0_elements(204) is a control-delay.
    cp_element_204_delay: control_delay_element  generic map(name => " 204_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(157), ack => testConfigure_CP_0_elements(204), clk => clk, reset =>reset);
    -- CP-element group 205:  transition  delay-element  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	164 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	170 
    -- CP-element group 205:  members (1) 
      -- CP-element group 205: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/ptr_deref_594_ptr_deref_624_delay
      -- 
    -- Element group testConfigure_CP_0_elements(205) is a control-delay.
    cp_element_205_delay: control_delay_element  generic map(name => " 205_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(164), ack => testConfigure_CP_0_elements(205), clk => clk, reset =>reset);
    -- CP-element group 206:  transition  delay-element  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	120 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	128 
    -- CP-element group 206:  members (1) 
      -- CP-element group 206: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/STORE_padding_452_STORE_padding_477_delay
      -- 
    -- Element group testConfigure_CP_0_elements(206) is a control-delay.
    cp_element_206_delay: control_delay_element  generic map(name => " 206_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(120), ack => testConfigure_CP_0_elements(206), clk => clk, reset =>reset);
    -- CP-element group 207:  branch  join  transition  place  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	121 
    -- CP-element group 207: 	130 
    -- CP-element group 207: 	137 
    -- CP-element group 207: 	144 
    -- CP-element group 207: 	151 
    -- CP-element group 207: 	158 
    -- CP-element group 207: 	165 
    -- CP-element group 207: 	172 
    -- CP-element group 207: 	176 
    -- CP-element group 207: 	180 
    -- CP-element group 207: 	184 
    -- CP-element group 207: 	188 
    -- CP-element group 207: 	192 
    -- CP-element group 207: 	196 
    -- CP-element group 207: 	200 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207: 	209 
    -- CP-element group 207:  members (10) 
      -- CP-element group 207: 	 branch_block_stmt_34/if_stmt_770_else_link/$entry
      -- CP-element group 207: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769__exit__
      -- CP-element group 207: 	 branch_block_stmt_34/if_stmt_770__entry__
      -- CP-element group 207: 	 branch_block_stmt_34/assign_stmt_454_to_assign_stmt_769/$exit
      -- CP-element group 207: 	 branch_block_stmt_34/R_cmp151299_771_place
      -- CP-element group 207: 	 branch_block_stmt_34/if_stmt_770_if_link/$entry
      -- CP-element group 207: 	 branch_block_stmt_34/if_stmt_770_eval_test/branch_req
      -- CP-element group 207: 	 branch_block_stmt_34/if_stmt_770_eval_test/$exit
      -- CP-element group 207: 	 branch_block_stmt_34/if_stmt_770_eval_test/$entry
      -- CP-element group 207: 	 branch_block_stmt_34/if_stmt_770_dead_link/$entry
      -- 
    branch_req_2363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(207), ack => if_stmt_770_branch_req_0); -- 
    testConfigure_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 14) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1);
      constant place_markings: IntegerArray(0 to 14)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0);
      constant place_delays: IntegerArray(0 to 14) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 15); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(121) & testConfigure_CP_0_elements(130) & testConfigure_CP_0_elements(137) & testConfigure_CP_0_elements(144) & testConfigure_CP_0_elements(151) & testConfigure_CP_0_elements(158) & testConfigure_CP_0_elements(165) & testConfigure_CP_0_elements(172) & testConfigure_CP_0_elements(176) & testConfigure_CP_0_elements(180) & testConfigure_CP_0_elements(184) & testConfigure_CP_0_elements(188) & testConfigure_CP_0_elements(192) & testConfigure_CP_0_elements(196) & testConfigure_CP_0_elements(200);
      gj_testConfigure_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 15, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	212 
    -- CP-element group 208: 	213 
    -- CP-element group 208:  members (18) 
      -- CP-element group 208: 	 branch_block_stmt_34/if_stmt_770_if_link/$exit
      -- CP-element group 208: 	 branch_block_stmt_34/if_stmt_770_if_link/if_choice_transition
      -- CP-element group 208: 	 branch_block_stmt_34/merge_stmt_791__exit__
      -- CP-element group 208: 	 branch_block_stmt_34/assign_stmt_797_to_assign_stmt_826__entry__
      -- CP-element group 208: 	 branch_block_stmt_34/assign_stmt_797_to_assign_stmt_826/type_cast_812_update_start_
      -- CP-element group 208: 	 branch_block_stmt_34/assign_stmt_797_to_assign_stmt_826/type_cast_812_sample_start_
      -- CP-element group 208: 	 branch_block_stmt_34/assign_stmt_797_to_assign_stmt_826/type_cast_812_Sample/$entry
      -- CP-element group 208: 	 branch_block_stmt_34/assign_stmt_797_to_assign_stmt_826/$entry
      -- CP-element group 208: 	 branch_block_stmt_34/forx_xend91_bbx_xnph301
      -- CP-element group 208: 	 branch_block_stmt_34/assign_stmt_797_to_assign_stmt_826/type_cast_812_Sample/rr
      -- CP-element group 208: 	 branch_block_stmt_34/assign_stmt_797_to_assign_stmt_826/type_cast_812_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_34/assign_stmt_797_to_assign_stmt_826/type_cast_812_Update/cr
      -- CP-element group 208: 	 branch_block_stmt_34/forx_xend91_bbx_xnph301_PhiReq/$entry
      -- CP-element group 208: 	 branch_block_stmt_34/forx_xend91_bbx_xnph301_PhiReq/$exit
      -- CP-element group 208: 	 branch_block_stmt_34/merge_stmt_791_PhiReqMerge
      -- CP-element group 208: 	 branch_block_stmt_34/merge_stmt_791_PhiAck/$entry
      -- CP-element group 208: 	 branch_block_stmt_34/merge_stmt_791_PhiAck/$exit
      -- CP-element group 208: 	 branch_block_stmt_34/merge_stmt_791_PhiAck/dummy
      -- 
    if_choice_transition_2368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_770_branch_ack_1, ack => testConfigure_CP_0_elements(208)); -- 
    rr_2407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(208), ack => type_cast_812_inst_req_0); -- 
    cr_2412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(208), ack => type_cast_812_inst_req_1); -- 
    -- CP-element group 209:  transition  place  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	387 
    -- CP-element group 209:  members (5) 
      -- CP-element group 209: 	 branch_block_stmt_34/if_stmt_770_else_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_34/forx_xend91_forx_xcond207x_xpreheader
      -- CP-element group 209: 	 branch_block_stmt_34/if_stmt_770_else_link/else_choice_transition
      -- CP-element group 209: 	 branch_block_stmt_34/forx_xend91_forx_xcond207x_xpreheader_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_34/forx_xend91_forx_xcond207x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_2372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_770_branch_ack_0, ack => testConfigure_CP_0_elements(209)); -- 
    -- CP-element group 210:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	387 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	256 
    -- CP-element group 210: 	257 
    -- CP-element group 210:  members (18) 
      -- CP-element group 210: 	 branch_block_stmt_34/merge_stmt_998__exit__
      -- CP-element group 210: 	 branch_block_stmt_34/assign_stmt_1004_to_assign_stmt_1033__entry__
      -- CP-element group 210: 	 branch_block_stmt_34/forx_xcond207x_xpreheader_bbx_xnph297
      -- CP-element group 210: 	 branch_block_stmt_34/if_stmt_785_if_link/if_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_34/if_stmt_785_if_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_34/assign_stmt_1004_to_assign_stmt_1033/$entry
      -- CP-element group 210: 	 branch_block_stmt_34/assign_stmt_1004_to_assign_stmt_1033/type_cast_1019_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_34/assign_stmt_1004_to_assign_stmt_1033/type_cast_1019_update_start_
      -- CP-element group 210: 	 branch_block_stmt_34/assign_stmt_1004_to_assign_stmt_1033/type_cast_1019_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_34/assign_stmt_1004_to_assign_stmt_1033/type_cast_1019_Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_34/assign_stmt_1004_to_assign_stmt_1033/type_cast_1019_Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_34/assign_stmt_1004_to_assign_stmt_1033/type_cast_1019_Update/cr
      -- CP-element group 210: 	 branch_block_stmt_34/forx_xcond207x_xpreheader_bbx_xnph297_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_34/forx_xcond207x_xpreheader_bbx_xnph297_PhiReq/$exit
      -- CP-element group 210: 	 branch_block_stmt_34/merge_stmt_998_PhiReqMerge
      -- CP-element group 210: 	 branch_block_stmt_34/merge_stmt_998_PhiAck/$entry
      -- CP-element group 210: 	 branch_block_stmt_34/merge_stmt_998_PhiAck/$exit
      -- CP-element group 210: 	 branch_block_stmt_34/merge_stmt_998_PhiAck/dummy
      -- 
    if_choice_transition_2390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_785_branch_ack_1, ack => testConfigure_CP_0_elements(210)); -- 
    rr_2766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(210), ack => type_cast_1019_inst_req_0); -- 
    cr_2771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(210), ack => type_cast_1019_inst_req_1); -- 
    -- CP-element group 211:  transition  place  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	387 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	400 
    -- CP-element group 211:  members (5) 
      -- CP-element group 211: 	 branch_block_stmt_34/forx_xcond207x_xpreheader_forx_xend267
      -- CP-element group 211: 	 branch_block_stmt_34/if_stmt_785_else_link/else_choice_transition
      -- CP-element group 211: 	 branch_block_stmt_34/if_stmt_785_else_link/$exit
      -- CP-element group 211: 	 branch_block_stmt_34/forx_xcond207x_xpreheader_forx_xend267_PhiReq/$entry
      -- CP-element group 211: 	 branch_block_stmt_34/forx_xcond207x_xpreheader_forx_xend267_PhiReq/$exit
      -- 
    else_choice_transition_2394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_785_branch_ack_0, ack => testConfigure_CP_0_elements(211)); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	208 
    -- CP-element group 212: successors 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_34/assign_stmt_797_to_assign_stmt_826/type_cast_812_sample_completed_
      -- CP-element group 212: 	 branch_block_stmt_34/assign_stmt_797_to_assign_stmt_826/type_cast_812_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_34/assign_stmt_797_to_assign_stmt_826/type_cast_812_Sample/ra
      -- 
    ra_2408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_812_inst_ack_0, ack => testConfigure_CP_0_elements(212)); -- 
    -- CP-element group 213:  transition  place  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	208 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	388 
    -- CP-element group 213:  members (9) 
      -- CP-element group 213: 	 branch_block_stmt_34/assign_stmt_797_to_assign_stmt_826/$exit
      -- CP-element group 213: 	 branch_block_stmt_34/assign_stmt_797_to_assign_stmt_826__exit__
      -- CP-element group 213: 	 branch_block_stmt_34/bbx_xnph301_forx_xbody153
      -- CP-element group 213: 	 branch_block_stmt_34/assign_stmt_797_to_assign_stmt_826/type_cast_812_update_completed_
      -- CP-element group 213: 	 branch_block_stmt_34/assign_stmt_797_to_assign_stmt_826/type_cast_812_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_34/assign_stmt_797_to_assign_stmt_826/type_cast_812_Update/ca
      -- CP-element group 213: 	 branch_block_stmt_34/bbx_xnph301_forx_xbody153_PhiReq/$entry
      -- CP-element group 213: 	 branch_block_stmt_34/bbx_xnph301_forx_xbody153_PhiReq/phi_stmt_829/$entry
      -- CP-element group 213: 	 branch_block_stmt_34/bbx_xnph301_forx_xbody153_PhiReq/phi_stmt_829/phi_stmt_829_sources/$entry
      -- 
    ca_2413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_812_inst_ack_1, ack => testConfigure_CP_0_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	393 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	253 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_final_index_sum_regn_Sample/ack
      -- CP-element group 214: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_final_index_sum_regn_Sample/$exit
      -- CP-element group 214: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_final_index_sum_regn_sample_complete
      -- 
    ack_2442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_841_index_offset_ack_0, ack => testConfigure_CP_0_elements(214)); -- 
    -- CP-element group 215:  transition  input  output  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	393 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215:  members (11) 
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_final_index_sum_regn_Update/ack
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_final_index_sum_regn_Update/$exit
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_base_plus_offset/sum_rename_req
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_base_plus_offset/$exit
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/addr_of_842_sample_start_
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_base_plus_offset/$entry
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_root_address_calculated
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_offset_calculated
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/addr_of_842_request/req
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/addr_of_842_request/$entry
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_base_plus_offset/sum_rename_ack
      -- 
    ack_2447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_841_index_offset_ack_1, ack => testConfigure_CP_0_elements(215)); -- 
    req_2456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(215), ack => addr_of_842_final_reg_req_0); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/addr_of_842_sample_completed_
      -- CP-element group 216: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/addr_of_842_request/ack
      -- CP-element group 216: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/addr_of_842_request/$exit
      -- 
    ack_2457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_842_final_reg_ack_0, ack => testConfigure_CP_0_elements(216)); -- 
    -- CP-element group 217:  fork  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	393 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	250 
    -- CP-element group 217:  members (19) 
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/addr_of_842_update_completed_
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/addr_of_842_complete/ack
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/addr_of_842_complete/$exit
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_base_address_calculated
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_word_address_calculated
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_root_address_calculated
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_base_address_resized
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_base_addr_resize/$entry
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_base_addr_resize/$exit
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_base_addr_resize/base_resize_req
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_base_addr_resize/base_resize_ack
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_base_plus_offset/$entry
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_base_plus_offset/$exit
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_base_plus_offset/sum_rename_req
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_base_plus_offset/sum_rename_ack
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_word_addrgen/$entry
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_word_addrgen/$exit
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_word_addrgen/root_register_req
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_word_addrgen/root_register_ack
      -- 
    ack_2462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_842_final_reg_ack_1, ack => testConfigure_CP_0_elements(217)); -- 
    -- CP-element group 218:  transition  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	393 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (6) 
      -- CP-element group 218: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_845_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_845_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_845_Sample/ra
      -- CP-element group 218: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_845_Sample/$exit
      -- CP-element group 218: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_845_update_start_
      -- CP-element group 218: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_845_sample_completed_
      -- 
    ra_2471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_845_inst_ack_0, ack => testConfigure_CP_0_elements(218)); -- 
    cr_2475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(218), ack => RPIPE_ConvTranspose_input_pipe_845_inst_req_1); -- 
    -- CP-element group 219:  fork  transition  input  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	220 
    -- CP-element group 219: 	222 
    -- CP-element group 219:  members (9) 
      -- CP-element group 219: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_845_Update/ca
      -- CP-element group 219: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_849_sample_start_
      -- CP-element group 219: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_845_Update/$exit
      -- CP-element group 219: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_849_Sample/$entry
      -- CP-element group 219: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_845_update_completed_
      -- CP-element group 219: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_858_Sample/rr
      -- CP-element group 219: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_858_Sample/$entry
      -- CP-element group 219: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_858_sample_start_
      -- CP-element group 219: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_849_Sample/rr
      -- 
    ca_2476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_845_inst_ack_1, ack => testConfigure_CP_0_elements(219)); -- 
    rr_2484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(219), ack => type_cast_849_inst_req_0); -- 
    rr_2498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(219), ack => RPIPE_ConvTranspose_input_pipe_858_inst_req_0); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	219 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_849_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_849_Sample/ra
      -- CP-element group 220: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_849_Sample/$exit
      -- 
    ra_2485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_849_inst_ack_0, ack => testConfigure_CP_0_elements(220)); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	393 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	250 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_849_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_849_Update/ca
      -- CP-element group 221: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_849_Update/$exit
      -- 
    ca_2490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_849_inst_ack_1, ack => testConfigure_CP_0_elements(221)); -- 
    -- CP-element group 222:  transition  input  output  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	219 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (6) 
      -- CP-element group 222: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_858_Update/cr
      -- CP-element group 222: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_858_Update/$entry
      -- CP-element group 222: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_858_Sample/ra
      -- CP-element group 222: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_858_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_858_update_start_
      -- CP-element group 222: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_858_sample_completed_
      -- 
    ra_2499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_858_inst_ack_0, ack => testConfigure_CP_0_elements(222)); -- 
    cr_2503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(222), ack => RPIPE_ConvTranspose_input_pipe_858_inst_req_1); -- 
    -- CP-element group 223:  fork  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223: 	226 
    -- CP-element group 223:  members (9) 
      -- CP-element group 223: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_862_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_862_Sample/$entry
      -- CP-element group 223: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_862_Sample/rr
      -- CP-element group 223: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_876_Sample/$entry
      -- CP-element group 223: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_858_Update/ca
      -- CP-element group 223: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_858_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_876_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_858_update_completed_
      -- CP-element group 223: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_876_Sample/rr
      -- 
    ca_2504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_858_inst_ack_1, ack => testConfigure_CP_0_elements(223)); -- 
    rr_2512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(223), ack => type_cast_862_inst_req_0); -- 
    rr_2526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(223), ack => RPIPE_ConvTranspose_input_pipe_876_inst_req_0); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_862_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_862_Sample/$exit
      -- CP-element group 224: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_862_Sample/ra
      -- 
    ra_2513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_862_inst_ack_0, ack => testConfigure_CP_0_elements(224)); -- 
    -- CP-element group 225:  transition  input  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	393 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	250 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_862_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_862_Update/$exit
      -- CP-element group 225: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_862_Update/ca
      -- 
    ca_2518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_862_inst_ack_1, ack => testConfigure_CP_0_elements(225)); -- 
    -- CP-element group 226:  transition  input  output  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	223 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	227 
    -- CP-element group 226:  members (6) 
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_876_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_876_Update/cr
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_876_Update/$entry
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_876_update_start_
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_876_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_876_Sample/ra
      -- 
    ra_2527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_876_inst_ack_0, ack => testConfigure_CP_0_elements(226)); -- 
    cr_2531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(226), ack => RPIPE_ConvTranspose_input_pipe_876_inst_req_1); -- 
    -- CP-element group 227:  fork  transition  input  output  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	226 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227: 	230 
    -- CP-element group 227:  members (9) 
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_880_Sample/$entry
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_876_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_876_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_880_Sample/rr
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_876_Update/ca
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_894_Sample/rr
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_894_Sample/$entry
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_880_sample_start_
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_894_sample_start_
      -- 
    ca_2532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_876_inst_ack_1, ack => testConfigure_CP_0_elements(227)); -- 
    rr_2540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(227), ack => type_cast_880_inst_req_0); -- 
    rr_2554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(227), ack => RPIPE_ConvTranspose_input_pipe_894_inst_req_0); -- 
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_880_Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_880_Sample/ra
      -- CP-element group 228: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_880_sample_completed_
      -- 
    ra_2541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_880_inst_ack_0, ack => testConfigure_CP_0_elements(228)); -- 
    -- CP-element group 229:  transition  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	393 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	250 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_880_Update/ca
      -- CP-element group 229: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_880_update_completed_
      -- CP-element group 229: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_880_Update/$exit
      -- 
    ca_2546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_880_inst_ack_1, ack => testConfigure_CP_0_elements(229)); -- 
    -- CP-element group 230:  transition  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	227 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	231 
    -- CP-element group 230:  members (6) 
      -- CP-element group 230: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_894_Update/cr
      -- CP-element group 230: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_894_Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_894_Sample/ra
      -- CP-element group 230: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_894_Sample/$exit
      -- CP-element group 230: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_894_update_start_
      -- CP-element group 230: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_894_sample_completed_
      -- 
    ra_2555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_894_inst_ack_0, ack => testConfigure_CP_0_elements(230)); -- 
    cr_2559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(230), ack => RPIPE_ConvTranspose_input_pipe_894_inst_req_1); -- 
    -- CP-element group 231:  fork  transition  input  output  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231: 	234 
    -- CP-element group 231:  members (9) 
      -- CP-element group 231: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_898_sample_start_
      -- CP-element group 231: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_912_sample_start_
      -- CP-element group 231: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_894_Update/ca
      -- CP-element group 231: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_894_Update/$exit
      -- CP-element group 231: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_912_Sample/rr
      -- CP-element group 231: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_894_update_completed_
      -- CP-element group 231: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_898_Sample/rr
      -- CP-element group 231: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_898_Sample/$entry
      -- CP-element group 231: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_912_Sample/$entry
      -- 
    ca_2560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_894_inst_ack_1, ack => testConfigure_CP_0_elements(231)); -- 
    rr_2568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(231), ack => type_cast_898_inst_req_0); -- 
    rr_2582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(231), ack => RPIPE_ConvTranspose_input_pipe_912_inst_req_0); -- 
    -- CP-element group 232:  transition  input  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_898_sample_completed_
      -- CP-element group 232: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_898_Sample/ra
      -- CP-element group 232: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_898_Sample/$exit
      -- 
    ra_2569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_898_inst_ack_0, ack => testConfigure_CP_0_elements(232)); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	393 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	250 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_898_update_completed_
      -- CP-element group 233: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_898_Update/ca
      -- CP-element group 233: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_898_Update/$exit
      -- 
    ca_2574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_898_inst_ack_1, ack => testConfigure_CP_0_elements(233)); -- 
    -- CP-element group 234:  transition  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	231 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234:  members (6) 
      -- CP-element group 234: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_912_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_912_sample_completed_
      -- CP-element group 234: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_912_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_912_Sample/ra
      -- CP-element group 234: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_912_Sample/$exit
      -- CP-element group 234: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_912_update_start_
      -- 
    ra_2583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_912_inst_ack_0, ack => testConfigure_CP_0_elements(234)); -- 
    cr_2587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(234), ack => RPIPE_ConvTranspose_input_pipe_912_inst_req_1); -- 
    -- CP-element group 235:  fork  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235: 	238 
    -- CP-element group 235:  members (9) 
      -- CP-element group 235: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_912_Update/$exit
      -- CP-element group 235: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_916_Sample/rr
      -- CP-element group 235: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_916_Sample/$entry
      -- CP-element group 235: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_916_sample_start_
      -- CP-element group 235: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_912_update_completed_
      -- CP-element group 235: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_912_Update/ca
      -- CP-element group 235: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_930_sample_start_
      -- CP-element group 235: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_930_Sample/$entry
      -- CP-element group 235: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_930_Sample/rr
      -- 
    ca_2588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_912_inst_ack_1, ack => testConfigure_CP_0_elements(235)); -- 
    rr_2596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(235), ack => type_cast_916_inst_req_0); -- 
    rr_2610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(235), ack => RPIPE_ConvTranspose_input_pipe_930_inst_req_0); -- 
    -- CP-element group 236:  transition  input  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_916_sample_completed_
      -- CP-element group 236: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_916_Sample/ra
      -- CP-element group 236: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_916_Sample/$exit
      -- 
    ra_2597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_916_inst_ack_0, ack => testConfigure_CP_0_elements(236)); -- 
    -- CP-element group 237:  transition  input  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	393 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	250 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_916_Update/ca
      -- CP-element group 237: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_916_Update/$exit
      -- CP-element group 237: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_916_update_completed_
      -- 
    ca_2602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_916_inst_ack_1, ack => testConfigure_CP_0_elements(237)); -- 
    -- CP-element group 238:  transition  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	235 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_930_sample_completed_
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_930_update_start_
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_930_Sample/$exit
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_930_Sample/ra
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_930_Update/$entry
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_930_Update/cr
      -- 
    ra_2611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_930_inst_ack_0, ack => testConfigure_CP_0_elements(238)); -- 
    cr_2615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(238), ack => RPIPE_ConvTranspose_input_pipe_930_inst_req_1); -- 
    -- CP-element group 239:  fork  transition  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239: 	242 
    -- CP-element group 239:  members (9) 
      -- CP-element group 239: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_930_update_completed_
      -- CP-element group 239: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_930_Update/$exit
      -- CP-element group 239: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_930_Update/ca
      -- CP-element group 239: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_934_sample_start_
      -- CP-element group 239: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_934_Sample/$entry
      -- CP-element group 239: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_934_Sample/rr
      -- CP-element group 239: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_948_sample_start_
      -- CP-element group 239: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_948_Sample/$entry
      -- CP-element group 239: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_948_Sample/rr
      -- 
    ca_2616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_930_inst_ack_1, ack => testConfigure_CP_0_elements(239)); -- 
    rr_2624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(239), ack => type_cast_934_inst_req_0); -- 
    rr_2638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(239), ack => RPIPE_ConvTranspose_input_pipe_948_inst_req_0); -- 
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_934_sample_completed_
      -- CP-element group 240: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_934_Sample/$exit
      -- CP-element group 240: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_934_Sample/ra
      -- 
    ra_2625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_934_inst_ack_0, ack => testConfigure_CP_0_elements(240)); -- 
    -- CP-element group 241:  transition  input  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	393 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	250 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_934_update_completed_
      -- CP-element group 241: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_934_Update/$exit
      -- CP-element group 241: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_934_Update/ca
      -- 
    ca_2630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_934_inst_ack_1, ack => testConfigure_CP_0_elements(241)); -- 
    -- CP-element group 242:  transition  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	239 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (6) 
      -- CP-element group 242: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_948_sample_completed_
      -- CP-element group 242: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_948_update_start_
      -- CP-element group 242: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_948_Sample/$exit
      -- CP-element group 242: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_948_Sample/ra
      -- CP-element group 242: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_948_Update/$entry
      -- CP-element group 242: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_948_Update/cr
      -- 
    ra_2639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_948_inst_ack_0, ack => testConfigure_CP_0_elements(242)); -- 
    cr_2643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(242), ack => RPIPE_ConvTranspose_input_pipe_948_inst_req_1); -- 
    -- CP-element group 243:  fork  transition  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243: 	246 
    -- CP-element group 243:  members (9) 
      -- CP-element group 243: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_948_update_completed_
      -- CP-element group 243: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_948_Update/$exit
      -- CP-element group 243: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_948_Update/ca
      -- CP-element group 243: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_952_sample_start_
      -- CP-element group 243: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_952_Sample/$entry
      -- CP-element group 243: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_952_Sample/rr
      -- CP-element group 243: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_966_sample_start_
      -- CP-element group 243: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_966_Sample/$entry
      -- CP-element group 243: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_966_Sample/rr
      -- 
    ca_2644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_948_inst_ack_1, ack => testConfigure_CP_0_elements(243)); -- 
    rr_2652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(243), ack => type_cast_952_inst_req_0); -- 
    rr_2666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(243), ack => RPIPE_ConvTranspose_input_pipe_966_inst_req_0); -- 
    -- CP-element group 244:  transition  input  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_952_sample_completed_
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_952_Sample/$exit
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_952_Sample/ra
      -- 
    ra_2653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_952_inst_ack_0, ack => testConfigure_CP_0_elements(244)); -- 
    -- CP-element group 245:  transition  input  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	393 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	250 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_952_update_completed_
      -- CP-element group 245: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_952_Update/$exit
      -- CP-element group 245: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_952_Update/ca
      -- 
    ca_2658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_952_inst_ack_1, ack => testConfigure_CP_0_elements(245)); -- 
    -- CP-element group 246:  transition  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	243 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (6) 
      -- CP-element group 246: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_966_sample_completed_
      -- CP-element group 246: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_966_update_start_
      -- CP-element group 246: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_966_Sample/$exit
      -- CP-element group 246: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_966_Sample/ra
      -- CP-element group 246: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_966_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_966_Update/cr
      -- 
    ra_2667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_966_inst_ack_0, ack => testConfigure_CP_0_elements(246)); -- 
    cr_2671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(246), ack => RPIPE_ConvTranspose_input_pipe_966_inst_req_1); -- 
    -- CP-element group 247:  transition  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_966_update_completed_
      -- CP-element group 247: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_966_Update/$exit
      -- CP-element group 247: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_966_Update/ca
      -- CP-element group 247: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_970_sample_start_
      -- CP-element group 247: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_970_Sample/$entry
      -- CP-element group 247: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_970_Sample/rr
      -- 
    ca_2672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_966_inst_ack_1, ack => testConfigure_CP_0_elements(247)); -- 
    rr_2680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(247), ack => type_cast_970_inst_req_0); -- 
    -- CP-element group 248:  transition  input  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_970_sample_completed_
      -- CP-element group 248: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_970_Sample/$exit
      -- CP-element group 248: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_970_Sample/ra
      -- 
    ra_2681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_970_inst_ack_0, ack => testConfigure_CP_0_elements(248)); -- 
    -- CP-element group 249:  transition  input  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	393 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_970_update_completed_
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_970_Update/$exit
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_970_Update/ca
      -- 
    ca_2686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_970_inst_ack_1, ack => testConfigure_CP_0_elements(249)); -- 
    -- CP-element group 250:  join  transition  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	217 
    -- CP-element group 250: 	221 
    -- CP-element group 250: 	225 
    -- CP-element group 250: 	229 
    -- CP-element group 250: 	233 
    -- CP-element group 250: 	237 
    -- CP-element group 250: 	241 
    -- CP-element group 250: 	245 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (9) 
      -- CP-element group 250: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_Sample/ptr_deref_978_Split/$entry
      -- CP-element group 250: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_Sample/ptr_deref_978_Split/$exit
      -- CP-element group 250: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_Sample/ptr_deref_978_Split/split_req
      -- CP-element group 250: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_Sample/ptr_deref_978_Split/split_ack
      -- CP-element group 250: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_Sample/word_access_start/$entry
      -- CP-element group 250: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_Sample/word_access_start/word_0/$entry
      -- CP-element group 250: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_Sample/word_access_start/word_0/rr
      -- 
    rr_2724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(250), ack => ptr_deref_978_store_0_req_0); -- 
    testConfigure_cp_element_group_250: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_250"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(217) & testConfigure_CP_0_elements(221) & testConfigure_CP_0_elements(225) & testConfigure_CP_0_elements(229) & testConfigure_CP_0_elements(233) & testConfigure_CP_0_elements(237) & testConfigure_CP_0_elements(241) & testConfigure_CP_0_elements(245) & testConfigure_CP_0_elements(249);
      gj_testConfigure_cp_element_group_250 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(250), clk => clk, reset => reset); --
    end block;
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251:  members (5) 
      -- CP-element group 251: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_Sample/word_access_start/$exit
      -- CP-element group 251: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_Sample/word_access_start/word_0/$exit
      -- CP-element group 251: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_Sample/word_access_start/word_0/ra
      -- 
    ra_2725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_978_store_0_ack_0, ack => testConfigure_CP_0_elements(251)); -- 
    -- CP-element group 252:  transition  input  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	393 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (5) 
      -- CP-element group 252: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_Update/word_access_complete/$exit
      -- CP-element group 252: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_Update/word_access_complete/word_0/$exit
      -- CP-element group 252: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_Update/word_access_complete/word_0/ca
      -- 
    ca_2736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_978_store_0_ack_1, ack => testConfigure_CP_0_elements(252)); -- 
    -- CP-element group 253:  branch  join  transition  place  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	214 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (10) 
      -- CP-element group 253: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991__exit__
      -- CP-element group 253: 	 branch_block_stmt_34/if_stmt_992__entry__
      -- CP-element group 253: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/$exit
      -- CP-element group 253: 	 branch_block_stmt_34/if_stmt_992_dead_link/$entry
      -- CP-element group 253: 	 branch_block_stmt_34/if_stmt_992_eval_test/$entry
      -- CP-element group 253: 	 branch_block_stmt_34/if_stmt_992_eval_test/$exit
      -- CP-element group 253: 	 branch_block_stmt_34/if_stmt_992_eval_test/branch_req
      -- CP-element group 253: 	 branch_block_stmt_34/R_exitcond6_993_place
      -- CP-element group 253: 	 branch_block_stmt_34/if_stmt_992_if_link/$entry
      -- CP-element group 253: 	 branch_block_stmt_34/if_stmt_992_else_link/$entry
      -- 
    branch_req_2744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(253), ack => if_stmt_992_branch_req_0); -- 
    testConfigure_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(214) & testConfigure_CP_0_elements(252);
      gj_testConfigure_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  merge  transition  place  input  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	387 
    -- CP-element group 254:  members (13) 
      -- CP-element group 254: 	 branch_block_stmt_34/merge_stmt_776__exit__
      -- CP-element group 254: 	 branch_block_stmt_34/forx_xcond207x_xpreheaderx_xloopexit_forx_xcond207x_xpreheader
      -- CP-element group 254: 	 branch_block_stmt_34/if_stmt_992_if_link/$exit
      -- CP-element group 254: 	 branch_block_stmt_34/if_stmt_992_if_link/if_choice_transition
      -- CP-element group 254: 	 branch_block_stmt_34/forx_xbody153_forx_xcond207x_xpreheaderx_xloopexit
      -- CP-element group 254: 	 branch_block_stmt_34/forx_xbody153_forx_xcond207x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 254: 	 branch_block_stmt_34/forx_xbody153_forx_xcond207x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 254: 	 branch_block_stmt_34/merge_stmt_776_PhiReqMerge
      -- CP-element group 254: 	 branch_block_stmt_34/merge_stmt_776_PhiAck/$entry
      -- CP-element group 254: 	 branch_block_stmt_34/merge_stmt_776_PhiAck/$exit
      -- CP-element group 254: 	 branch_block_stmt_34/merge_stmt_776_PhiAck/dummy
      -- CP-element group 254: 	 branch_block_stmt_34/forx_xcond207x_xpreheaderx_xloopexit_forx_xcond207x_xpreheader_PhiReq/$entry
      -- CP-element group 254: 	 branch_block_stmt_34/forx_xcond207x_xpreheaderx_xloopexit_forx_xcond207x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_2749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_992_branch_ack_1, ack => testConfigure_CP_0_elements(254)); -- 
    -- CP-element group 255:  fork  transition  place  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	389 
    -- CP-element group 255: 	390 
    -- CP-element group 255:  members (12) 
      -- CP-element group 255: 	 branch_block_stmt_34/if_stmt_992_else_link/$exit
      -- CP-element group 255: 	 branch_block_stmt_34/if_stmt_992_else_link/else_choice_transition
      -- CP-element group 255: 	 branch_block_stmt_34/forx_xbody153_forx_xbody153
      -- CP-element group 255: 	 branch_block_stmt_34/forx_xbody153_forx_xbody153_PhiReq/$entry
      -- CP-element group 255: 	 branch_block_stmt_34/forx_xbody153_forx_xbody153_PhiReq/phi_stmt_829/$entry
      -- CP-element group 255: 	 branch_block_stmt_34/forx_xbody153_forx_xbody153_PhiReq/phi_stmt_829/phi_stmt_829_sources/$entry
      -- CP-element group 255: 	 branch_block_stmt_34/forx_xbody153_forx_xbody153_PhiReq/phi_stmt_829/phi_stmt_829_sources/type_cast_835/$entry
      -- CP-element group 255: 	 branch_block_stmt_34/forx_xbody153_forx_xbody153_PhiReq/phi_stmt_829/phi_stmt_829_sources/type_cast_835/SplitProtocol/$entry
      -- CP-element group 255: 	 branch_block_stmt_34/forx_xbody153_forx_xbody153_PhiReq/phi_stmt_829/phi_stmt_829_sources/type_cast_835/SplitProtocol/Sample/$entry
      -- CP-element group 255: 	 branch_block_stmt_34/forx_xbody153_forx_xbody153_PhiReq/phi_stmt_829/phi_stmt_829_sources/type_cast_835/SplitProtocol/Sample/rr
      -- CP-element group 255: 	 branch_block_stmt_34/forx_xbody153_forx_xbody153_PhiReq/phi_stmt_829/phi_stmt_829_sources/type_cast_835/SplitProtocol/Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_34/forx_xbody153_forx_xbody153_PhiReq/phi_stmt_829/phi_stmt_829_sources/type_cast_835/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_992_branch_ack_0, ack => testConfigure_CP_0_elements(255)); -- 
    rr_3949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(255), ack => type_cast_835_inst_req_0); -- 
    cr_3954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(255), ack => type_cast_835_inst_req_1); -- 
    -- CP-element group 256:  transition  input  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	210 
    -- CP-element group 256: successors 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_34/assign_stmt_1004_to_assign_stmt_1033/type_cast_1019_sample_completed_
      -- CP-element group 256: 	 branch_block_stmt_34/assign_stmt_1004_to_assign_stmt_1033/type_cast_1019_Sample/$exit
      -- CP-element group 256: 	 branch_block_stmt_34/assign_stmt_1004_to_assign_stmt_1033/type_cast_1019_Sample/ra
      -- 
    ra_2767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1019_inst_ack_0, ack => testConfigure_CP_0_elements(256)); -- 
    -- CP-element group 257:  transition  place  input  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	210 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	394 
    -- CP-element group 257:  members (9) 
      -- CP-element group 257: 	 branch_block_stmt_34/assign_stmt_1004_to_assign_stmt_1033__exit__
      -- CP-element group 257: 	 branch_block_stmt_34/bbx_xnph297_forx_xbody213
      -- CP-element group 257: 	 branch_block_stmt_34/assign_stmt_1004_to_assign_stmt_1033/$exit
      -- CP-element group 257: 	 branch_block_stmt_34/assign_stmt_1004_to_assign_stmt_1033/type_cast_1019_update_completed_
      -- CP-element group 257: 	 branch_block_stmt_34/assign_stmt_1004_to_assign_stmt_1033/type_cast_1019_Update/$exit
      -- CP-element group 257: 	 branch_block_stmt_34/assign_stmt_1004_to_assign_stmt_1033/type_cast_1019_Update/ca
      -- CP-element group 257: 	 branch_block_stmt_34/bbx_xnph297_forx_xbody213_PhiReq/$entry
      -- CP-element group 257: 	 branch_block_stmt_34/bbx_xnph297_forx_xbody213_PhiReq/phi_stmt_1036/$entry
      -- CP-element group 257: 	 branch_block_stmt_34/bbx_xnph297_forx_xbody213_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/$entry
      -- 
    ca_2772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1019_inst_ack_1, ack => testConfigure_CP_0_elements(257)); -- 
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	399 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	297 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_final_index_sum_regn_sample_complete
      -- CP-element group 258: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_final_index_sum_regn_Sample/$exit
      -- CP-element group 258: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_final_index_sum_regn_Sample/ack
      -- 
    ack_2801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1048_index_offset_ack_0, ack => testConfigure_CP_0_elements(258)); -- 
    -- CP-element group 259:  transition  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	399 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (11) 
      -- CP-element group 259: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/addr_of_1049_sample_start_
      -- CP-element group 259: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_root_address_calculated
      -- CP-element group 259: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_offset_calculated
      -- CP-element group 259: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_final_index_sum_regn_Update/$exit
      -- CP-element group 259: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_final_index_sum_regn_Update/ack
      -- CP-element group 259: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_base_plus_offset/$entry
      -- CP-element group 259: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_base_plus_offset/$exit
      -- CP-element group 259: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_base_plus_offset/sum_rename_req
      -- CP-element group 259: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_base_plus_offset/sum_rename_ack
      -- CP-element group 259: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/addr_of_1049_request/$entry
      -- CP-element group 259: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/addr_of_1049_request/req
      -- 
    ack_2806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1048_index_offset_ack_1, ack => testConfigure_CP_0_elements(259)); -- 
    req_2815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(259), ack => addr_of_1049_final_reg_req_0); -- 
    -- CP-element group 260:  transition  input  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/addr_of_1049_sample_completed_
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/addr_of_1049_request/$exit
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/addr_of_1049_request/ack
      -- 
    ack_2816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1049_final_reg_ack_0, ack => testConfigure_CP_0_elements(260)); -- 
    -- CP-element group 261:  fork  transition  input  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	399 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	294 
    -- CP-element group 261:  members (19) 
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/addr_of_1049_update_completed_
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/addr_of_1049_complete/$exit
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/addr_of_1049_complete/ack
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_base_address_calculated
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_word_address_calculated
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_root_address_calculated
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_base_address_resized
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_base_addr_resize/$entry
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_base_addr_resize/$exit
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_base_addr_resize/base_resize_req
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_base_addr_resize/base_resize_ack
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_base_plus_offset/$entry
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_base_plus_offset/$exit
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_base_plus_offset/sum_rename_req
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_base_plus_offset/sum_rename_ack
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_word_addrgen/$entry
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_word_addrgen/$exit
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_word_addrgen/root_register_req
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_word_addrgen/root_register_ack
      -- 
    ack_2821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1049_final_reg_ack_1, ack => testConfigure_CP_0_elements(261)); -- 
    -- CP-element group 262:  transition  input  output  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	399 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	263 
    -- CP-element group 262:  members (6) 
      -- CP-element group 262: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1052_sample_completed_
      -- CP-element group 262: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1052_update_start_
      -- CP-element group 262: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1052_Sample/$exit
      -- CP-element group 262: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1052_Sample/ra
      -- CP-element group 262: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1052_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1052_Update/cr
      -- 
    ra_2830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1052_inst_ack_0, ack => testConfigure_CP_0_elements(262)); -- 
    cr_2834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(262), ack => RPIPE_ConvTranspose_input_pipe_1052_inst_req_1); -- 
    -- CP-element group 263:  fork  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	262 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263: 	266 
    -- CP-element group 263:  members (9) 
      -- CP-element group 263: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1052_update_completed_
      -- CP-element group 263: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1052_Update/$exit
      -- CP-element group 263: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1052_Update/ca
      -- CP-element group 263: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1056_sample_start_
      -- CP-element group 263: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1056_Sample/$entry
      -- CP-element group 263: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1056_Sample/rr
      -- CP-element group 263: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1065_sample_start_
      -- CP-element group 263: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1065_Sample/$entry
      -- CP-element group 263: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1065_Sample/rr
      -- 
    ca_2835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1052_inst_ack_1, ack => testConfigure_CP_0_elements(263)); -- 
    rr_2843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(263), ack => type_cast_1056_inst_req_0); -- 
    rr_2857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(263), ack => RPIPE_ConvTranspose_input_pipe_1065_inst_req_0); -- 
    -- CP-element group 264:  transition  input  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1056_sample_completed_
      -- CP-element group 264: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1056_Sample/$exit
      -- CP-element group 264: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1056_Sample/ra
      -- 
    ra_2844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1056_inst_ack_0, ack => testConfigure_CP_0_elements(264)); -- 
    -- CP-element group 265:  transition  input  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	399 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	294 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1056_update_completed_
      -- CP-element group 265: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1056_Update/$exit
      -- CP-element group 265: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1056_Update/ca
      -- 
    ca_2849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1056_inst_ack_1, ack => testConfigure_CP_0_elements(265)); -- 
    -- CP-element group 266:  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	263 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (6) 
      -- CP-element group 266: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1065_sample_completed_
      -- CP-element group 266: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1065_update_start_
      -- CP-element group 266: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1065_Sample/$exit
      -- CP-element group 266: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1065_Sample/ra
      -- CP-element group 266: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1065_Update/$entry
      -- CP-element group 266: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1065_Update/cr
      -- 
    ra_2858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1065_inst_ack_0, ack => testConfigure_CP_0_elements(266)); -- 
    cr_2862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(266), ack => RPIPE_ConvTranspose_input_pipe_1065_inst_req_1); -- 
    -- CP-element group 267:  fork  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267: 	270 
    -- CP-element group 267:  members (9) 
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1065_update_completed_
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1065_Update/$exit
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1065_Update/ca
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1069_sample_start_
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1069_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1069_Sample/rr
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1083_sample_start_
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1083_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1083_Sample/rr
      -- 
    ca_2863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1065_inst_ack_1, ack => testConfigure_CP_0_elements(267)); -- 
    rr_2871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => type_cast_1069_inst_req_0); -- 
    rr_2885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => RPIPE_ConvTranspose_input_pipe_1083_inst_req_0); -- 
    -- CP-element group 268:  transition  input  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1069_sample_completed_
      -- CP-element group 268: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1069_Sample/$exit
      -- CP-element group 268: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1069_Sample/ra
      -- 
    ra_2872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1069_inst_ack_0, ack => testConfigure_CP_0_elements(268)); -- 
    -- CP-element group 269:  transition  input  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	399 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	294 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1069_update_completed_
      -- CP-element group 269: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1069_Update/$exit
      -- CP-element group 269: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1069_Update/ca
      -- 
    ca_2877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1069_inst_ack_1, ack => testConfigure_CP_0_elements(269)); -- 
    -- CP-element group 270:  transition  input  output  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	267 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (6) 
      -- CP-element group 270: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1083_sample_completed_
      -- CP-element group 270: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1083_update_start_
      -- CP-element group 270: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1083_Sample/$exit
      -- CP-element group 270: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1083_Sample/ra
      -- CP-element group 270: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1083_Update/$entry
      -- CP-element group 270: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1083_Update/cr
      -- 
    ra_2886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1083_inst_ack_0, ack => testConfigure_CP_0_elements(270)); -- 
    cr_2890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(270), ack => RPIPE_ConvTranspose_input_pipe_1083_inst_req_1); -- 
    -- CP-element group 271:  fork  transition  input  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271: 	274 
    -- CP-element group 271:  members (9) 
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1083_update_completed_
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1083_Update/$exit
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1083_Update/ca
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1087_sample_start_
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1087_Sample/$entry
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1087_Sample/rr
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1101_sample_start_
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1101_Sample/$entry
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1101_Sample/rr
      -- 
    ca_2891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1083_inst_ack_1, ack => testConfigure_CP_0_elements(271)); -- 
    rr_2899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(271), ack => type_cast_1087_inst_req_0); -- 
    rr_2913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(271), ack => RPIPE_ConvTranspose_input_pipe_1101_inst_req_0); -- 
    -- CP-element group 272:  transition  input  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1087_sample_completed_
      -- CP-element group 272: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1087_Sample/$exit
      -- CP-element group 272: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1087_Sample/ra
      -- 
    ra_2900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1087_inst_ack_0, ack => testConfigure_CP_0_elements(272)); -- 
    -- CP-element group 273:  transition  input  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	399 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	294 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1087_update_completed_
      -- CP-element group 273: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1087_Update/$exit
      -- CP-element group 273: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1087_Update/ca
      -- 
    ca_2905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1087_inst_ack_1, ack => testConfigure_CP_0_elements(273)); -- 
    -- CP-element group 274:  transition  input  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	271 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (6) 
      -- CP-element group 274: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1101_sample_completed_
      -- CP-element group 274: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1101_update_start_
      -- CP-element group 274: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1101_Sample/$exit
      -- CP-element group 274: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1101_Sample/ra
      -- CP-element group 274: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1101_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1101_Update/cr
      -- 
    ra_2914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1101_inst_ack_0, ack => testConfigure_CP_0_elements(274)); -- 
    cr_2918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(274), ack => RPIPE_ConvTranspose_input_pipe_1101_inst_req_1); -- 
    -- CP-element group 275:  fork  transition  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275: 	278 
    -- CP-element group 275:  members (9) 
      -- CP-element group 275: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1101_update_completed_
      -- CP-element group 275: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1101_Update/$exit
      -- CP-element group 275: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1101_Update/ca
      -- CP-element group 275: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1105_sample_start_
      -- CP-element group 275: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1105_Sample/$entry
      -- CP-element group 275: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1105_Sample/rr
      -- CP-element group 275: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1119_sample_start_
      -- CP-element group 275: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1119_Sample/$entry
      -- CP-element group 275: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1119_Sample/rr
      -- 
    ca_2919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1101_inst_ack_1, ack => testConfigure_CP_0_elements(275)); -- 
    rr_2927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(275), ack => type_cast_1105_inst_req_0); -- 
    rr_2941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(275), ack => RPIPE_ConvTranspose_input_pipe_1119_inst_req_0); -- 
    -- CP-element group 276:  transition  input  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1105_sample_completed_
      -- CP-element group 276: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1105_Sample/$exit
      -- CP-element group 276: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1105_Sample/ra
      -- 
    ra_2928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1105_inst_ack_0, ack => testConfigure_CP_0_elements(276)); -- 
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	399 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	294 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1105_update_completed_
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1105_Update/$exit
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1105_Update/ca
      -- 
    ca_2933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1105_inst_ack_1, ack => testConfigure_CP_0_elements(277)); -- 
    -- CP-element group 278:  transition  input  output  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	275 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (6) 
      -- CP-element group 278: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1119_sample_completed_
      -- CP-element group 278: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1119_update_start_
      -- CP-element group 278: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1119_Sample/$exit
      -- CP-element group 278: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1119_Sample/ra
      -- CP-element group 278: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1119_Update/$entry
      -- CP-element group 278: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1119_Update/cr
      -- 
    ra_2942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1119_inst_ack_0, ack => testConfigure_CP_0_elements(278)); -- 
    cr_2946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(278), ack => RPIPE_ConvTranspose_input_pipe_1119_inst_req_1); -- 
    -- CP-element group 279:  fork  transition  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279: 	282 
    -- CP-element group 279:  members (9) 
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1119_update_completed_
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1119_Update/$exit
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1119_Update/ca
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1123_sample_start_
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1123_Sample/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1123_Sample/rr
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1137_sample_start_
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1137_Sample/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1137_Sample/rr
      -- 
    ca_2947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1119_inst_ack_1, ack => testConfigure_CP_0_elements(279)); -- 
    rr_2955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(279), ack => type_cast_1123_inst_req_0); -- 
    rr_2969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(279), ack => RPIPE_ConvTranspose_input_pipe_1137_inst_req_0); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1123_sample_completed_
      -- CP-element group 280: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1123_Sample/$exit
      -- CP-element group 280: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1123_Sample/ra
      -- 
    ra_2956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1123_inst_ack_0, ack => testConfigure_CP_0_elements(280)); -- 
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	399 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	294 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1123_update_completed_
      -- CP-element group 281: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1123_Update/$exit
      -- CP-element group 281: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1123_Update/ca
      -- 
    ca_2961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1123_inst_ack_1, ack => testConfigure_CP_0_elements(281)); -- 
    -- CP-element group 282:  transition  input  output  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	279 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (6) 
      -- CP-element group 282: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1137_sample_completed_
      -- CP-element group 282: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1137_update_start_
      -- CP-element group 282: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1137_Sample/$exit
      -- CP-element group 282: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1137_Sample/ra
      -- CP-element group 282: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1137_Update/$entry
      -- CP-element group 282: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1137_Update/cr
      -- 
    ra_2970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1137_inst_ack_0, ack => testConfigure_CP_0_elements(282)); -- 
    cr_2974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(282), ack => RPIPE_ConvTranspose_input_pipe_1137_inst_req_1); -- 
    -- CP-element group 283:  fork  transition  input  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283: 	286 
    -- CP-element group 283:  members (9) 
      -- CP-element group 283: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1137_update_completed_
      -- CP-element group 283: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1137_Update/$exit
      -- CP-element group 283: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1137_Update/ca
      -- CP-element group 283: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1141_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1141_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1141_Sample/rr
      -- CP-element group 283: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1155_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1155_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1155_Sample/rr
      -- 
    ca_2975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1137_inst_ack_1, ack => testConfigure_CP_0_elements(283)); -- 
    rr_2983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(283), ack => type_cast_1141_inst_req_0); -- 
    rr_2997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(283), ack => RPIPE_ConvTranspose_input_pipe_1155_inst_req_0); -- 
    -- CP-element group 284:  transition  input  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1141_sample_completed_
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1141_Sample/$exit
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1141_Sample/ra
      -- 
    ra_2984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1141_inst_ack_0, ack => testConfigure_CP_0_elements(284)); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	399 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	294 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1141_update_completed_
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1141_Update/$exit
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1141_Update/ca
      -- 
    ca_2989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1141_inst_ack_1, ack => testConfigure_CP_0_elements(285)); -- 
    -- CP-element group 286:  transition  input  output  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	283 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286:  members (6) 
      -- CP-element group 286: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1155_sample_completed_
      -- CP-element group 286: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1155_update_start_
      -- CP-element group 286: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1155_Sample/$exit
      -- CP-element group 286: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1155_Sample/ra
      -- CP-element group 286: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1155_Update/$entry
      -- CP-element group 286: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1155_Update/cr
      -- 
    ra_2998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1155_inst_ack_0, ack => testConfigure_CP_0_elements(286)); -- 
    cr_3002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(286), ack => RPIPE_ConvTranspose_input_pipe_1155_inst_req_1); -- 
    -- CP-element group 287:  fork  transition  input  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287: 	290 
    -- CP-element group 287:  members (9) 
      -- CP-element group 287: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1155_update_completed_
      -- CP-element group 287: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1155_Update/$exit
      -- CP-element group 287: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1155_Update/ca
      -- CP-element group 287: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1159_sample_start_
      -- CP-element group 287: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1159_Sample/$entry
      -- CP-element group 287: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1159_Sample/rr
      -- CP-element group 287: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1173_sample_start_
      -- CP-element group 287: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1173_Sample/$entry
      -- CP-element group 287: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1173_Sample/rr
      -- 
    ca_3003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1155_inst_ack_1, ack => testConfigure_CP_0_elements(287)); -- 
    rr_3011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(287), ack => type_cast_1159_inst_req_0); -- 
    rr_3025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(287), ack => RPIPE_ConvTranspose_input_pipe_1173_inst_req_0); -- 
    -- CP-element group 288:  transition  input  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1159_sample_completed_
      -- CP-element group 288: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1159_Sample/$exit
      -- CP-element group 288: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1159_Sample/ra
      -- 
    ra_3012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1159_inst_ack_0, ack => testConfigure_CP_0_elements(288)); -- 
    -- CP-element group 289:  transition  input  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	399 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	294 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1159_update_completed_
      -- CP-element group 289: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1159_Update/$exit
      -- CP-element group 289: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1159_Update/ca
      -- 
    ca_3017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1159_inst_ack_1, ack => testConfigure_CP_0_elements(289)); -- 
    -- CP-element group 290:  transition  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	287 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (6) 
      -- CP-element group 290: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1173_sample_completed_
      -- CP-element group 290: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1173_update_start_
      -- CP-element group 290: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1173_Sample/$exit
      -- CP-element group 290: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1173_Sample/ra
      -- CP-element group 290: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1173_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1173_Update/cr
      -- 
    ra_3026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1173_inst_ack_0, ack => testConfigure_CP_0_elements(290)); -- 
    cr_3030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(290), ack => RPIPE_ConvTranspose_input_pipe_1173_inst_req_1); -- 
    -- CP-element group 291:  transition  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1173_update_completed_
      -- CP-element group 291: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1173_Update/$exit
      -- CP-element group 291: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1173_Update/ca
      -- CP-element group 291: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1177_sample_start_
      -- CP-element group 291: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1177_Sample/$entry
      -- CP-element group 291: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1177_Sample/rr
      -- 
    ca_3031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_1173_inst_ack_1, ack => testConfigure_CP_0_elements(291)); -- 
    rr_3039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(291), ack => type_cast_1177_inst_req_0); -- 
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1177_sample_completed_
      -- CP-element group 292: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1177_Sample/$exit
      -- CP-element group 292: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1177_Sample/ra
      -- 
    ra_3040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1177_inst_ack_0, ack => testConfigure_CP_0_elements(292)); -- 
    -- CP-element group 293:  transition  input  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	399 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1177_update_completed_
      -- CP-element group 293: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1177_Update/$exit
      -- CP-element group 293: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1177_Update/ca
      -- 
    ca_3045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1177_inst_ack_1, ack => testConfigure_CP_0_elements(293)); -- 
    -- CP-element group 294:  join  transition  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	261 
    -- CP-element group 294: 	265 
    -- CP-element group 294: 	269 
    -- CP-element group 294: 	273 
    -- CP-element group 294: 	277 
    -- CP-element group 294: 	281 
    -- CP-element group 294: 	285 
    -- CP-element group 294: 	289 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (9) 
      -- CP-element group 294: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_sample_start_
      -- CP-element group 294: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_Sample/ptr_deref_1185_Split/$entry
      -- CP-element group 294: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_Sample/ptr_deref_1185_Split/$exit
      -- CP-element group 294: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_Sample/ptr_deref_1185_Split/split_req
      -- CP-element group 294: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_Sample/ptr_deref_1185_Split/split_ack
      -- CP-element group 294: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_Sample/word_access_start/$entry
      -- CP-element group 294: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_Sample/word_access_start/word_0/$entry
      -- CP-element group 294: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_Sample/word_access_start/word_0/rr
      -- 
    rr_3083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(294), ack => ptr_deref_1185_store_0_req_0); -- 
    testConfigure_cp_element_group_294: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_294"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(261) & testConfigure_CP_0_elements(265) & testConfigure_CP_0_elements(269) & testConfigure_CP_0_elements(273) & testConfigure_CP_0_elements(277) & testConfigure_CP_0_elements(281) & testConfigure_CP_0_elements(285) & testConfigure_CP_0_elements(289) & testConfigure_CP_0_elements(293);
      gj_testConfigure_cp_element_group_294 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(294), clk => clk, reset => reset); --
    end block;
    -- CP-element group 295:  transition  input  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295:  members (5) 
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_sample_completed_
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_Sample/word_access_start/$exit
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_Sample/word_access_start/word_0/$exit
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_Sample/word_access_start/word_0/ra
      -- 
    ra_3084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1185_store_0_ack_0, ack => testConfigure_CP_0_elements(295)); -- 
    -- CP-element group 296:  transition  input  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	399 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296:  members (5) 
      -- CP-element group 296: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_update_completed_
      -- CP-element group 296: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_Update/word_access_complete/$exit
      -- CP-element group 296: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_Update/word_access_complete/word_0/$exit
      -- CP-element group 296: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_Update/word_access_complete/word_0/ca
      -- 
    ca_3095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1185_store_0_ack_1, ack => testConfigure_CP_0_elements(296)); -- 
    -- CP-element group 297:  branch  join  transition  place  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	258 
    -- CP-element group 297: 	296 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297: 	299 
    -- CP-element group 297:  members (10) 
      -- CP-element group 297: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198__exit__
      -- CP-element group 297: 	 branch_block_stmt_34/if_stmt_1199__entry__
      -- CP-element group 297: 	 branch_block_stmt_34/if_stmt_1199_eval_test/$entry
      -- CP-element group 297: 	 branch_block_stmt_34/if_stmt_1199_eval_test/$exit
      -- CP-element group 297: 	 branch_block_stmt_34/if_stmt_1199_eval_test/branch_req
      -- CP-element group 297: 	 branch_block_stmt_34/if_stmt_1199_if_link/$entry
      -- CP-element group 297: 	 branch_block_stmt_34/if_stmt_1199_else_link/$entry
      -- CP-element group 297: 	 branch_block_stmt_34/if_stmt_1199_dead_link/$entry
      -- CP-element group 297: 	 branch_block_stmt_34/R_exitcond_1200_place
      -- CP-element group 297: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/$exit
      -- 
    branch_req_3103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(297), ack => if_stmt_1199_branch_req_0); -- 
    testConfigure_cp_element_group_297: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_297"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(258) & testConfigure_CP_0_elements(296);
      gj_testConfigure_cp_element_group_297 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(297), clk => clk, reset => reset); --
    end block;
    -- CP-element group 298:  merge  transition  place  input  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	400 
    -- CP-element group 298:  members (13) 
      -- CP-element group 298: 	 branch_block_stmt_34/merge_stmt_1205__exit__
      -- CP-element group 298: 	 branch_block_stmt_34/forx_xend267x_xloopexit_forx_xend267
      -- CP-element group 298: 	 branch_block_stmt_34/if_stmt_1199_if_link/$exit
      -- CP-element group 298: 	 branch_block_stmt_34/if_stmt_1199_if_link/if_choice_transition
      -- CP-element group 298: 	 branch_block_stmt_34/forx_xbody213_forx_xend267x_xloopexit
      -- CP-element group 298: 	 branch_block_stmt_34/forx_xbody213_forx_xend267x_xloopexit_PhiReq/$entry
      -- CP-element group 298: 	 branch_block_stmt_34/forx_xbody213_forx_xend267x_xloopexit_PhiReq/$exit
      -- CP-element group 298: 	 branch_block_stmt_34/merge_stmt_1205_PhiReqMerge
      -- CP-element group 298: 	 branch_block_stmt_34/merge_stmt_1205_PhiAck/$entry
      -- CP-element group 298: 	 branch_block_stmt_34/merge_stmt_1205_PhiAck/$exit
      -- CP-element group 298: 	 branch_block_stmt_34/merge_stmt_1205_PhiAck/dummy
      -- CP-element group 298: 	 branch_block_stmt_34/forx_xend267x_xloopexit_forx_xend267_PhiReq/$entry
      -- CP-element group 298: 	 branch_block_stmt_34/forx_xend267x_xloopexit_forx_xend267_PhiReq/$exit
      -- 
    if_choice_transition_3108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1199_branch_ack_1, ack => testConfigure_CP_0_elements(298)); -- 
    -- CP-element group 299:  fork  transition  place  input  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	297 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	395 
    -- CP-element group 299: 	396 
    -- CP-element group 299:  members (12) 
      -- CP-element group 299: 	 branch_block_stmt_34/forx_xbody213_forx_xbody213
      -- CP-element group 299: 	 branch_block_stmt_34/if_stmt_1199_else_link/else_choice_transition
      -- CP-element group 299: 	 branch_block_stmt_34/if_stmt_1199_else_link/$exit
      -- CP-element group 299: 	 branch_block_stmt_34/forx_xbody213_forx_xbody213_PhiReq/$entry
      -- CP-element group 299: 	 branch_block_stmt_34/forx_xbody213_forx_xbody213_PhiReq/phi_stmt_1036/$entry
      -- CP-element group 299: 	 branch_block_stmt_34/forx_xbody213_forx_xbody213_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/$entry
      -- CP-element group 299: 	 branch_block_stmt_34/forx_xbody213_forx_xbody213_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/$entry
      -- CP-element group 299: 	 branch_block_stmt_34/forx_xbody213_forx_xbody213_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/SplitProtocol/$entry
      -- CP-element group 299: 	 branch_block_stmt_34/forx_xbody213_forx_xbody213_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/SplitProtocol/Sample/$entry
      -- CP-element group 299: 	 branch_block_stmt_34/forx_xbody213_forx_xbody213_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/SplitProtocol/Sample/rr
      -- CP-element group 299: 	 branch_block_stmt_34/forx_xbody213_forx_xbody213_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/SplitProtocol/Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_34/forx_xbody213_forx_xbody213_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1199_branch_ack_0, ack => testConfigure_CP_0_elements(299)); -- 
    rr_4003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(299), ack => type_cast_1042_inst_req_0); -- 
    cr_4008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(299), ack => type_cast_1042_inst_req_1); -- 
    -- CP-element group 300:  transition  input  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	401 
    -- CP-element group 300: successors 
    -- CP-element group 300:  members (5) 
      -- CP-element group 300: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_sample_completed_
      -- CP-element group 300: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_Sample/word_access_start/word_0/ra
      -- CP-element group 300: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_Sample/word_access_start/word_0/$exit
      -- CP-element group 300: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_Sample/word_access_start/$exit
      -- CP-element group 300: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_Sample/$exit
      -- 
    ra_3151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1218_load_0_ack_0, ack => testConfigure_CP_0_elements(300)); -- 
    -- CP-element group 301:  transition  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	401 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (12) 
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1222_Sample/rr
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1222_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_Update/ptr_deref_1218_Merge/$exit
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_Update/ptr_deref_1218_Merge/merge_req
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1222_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_Update/ptr_deref_1218_Merge/merge_ack
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_Update/ptr_deref_1218_Merge/$entry
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_Update/word_access_complete/word_0/ca
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_Update/word_access_complete/word_0/$exit
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_update_completed_
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_Update/word_access_complete/$exit
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_Update/$exit
      -- 
    ca_3162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1218_load_0_ack_1, ack => testConfigure_CP_0_elements(301)); -- 
    rr_3175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_1222_inst_req_0); -- 
    -- CP-element group 302:  transition  input  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1222_Sample/$exit
      -- CP-element group 302: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1222_Sample/ra
      -- CP-element group 302: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1222_sample_completed_
      -- 
    ra_3176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1222_inst_ack_0, ack => testConfigure_CP_0_elements(302)); -- 
    -- CP-element group 303:  transition  input  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	401 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	312 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1222_Update/$exit
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1222_update_completed_
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1222_Update/ca
      -- 
    ca_3181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1222_inst_ack_1, ack => testConfigure_CP_0_elements(303)); -- 
    -- CP-element group 304:  transition  input  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	401 
    -- CP-element group 304: successors 
    -- CP-element group 304:  members (5) 
      -- CP-element group 304: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_sample_completed_
      -- CP-element group 304: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_Sample/word_access_start/word_0/ra
      -- CP-element group 304: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_Sample/word_access_start/word_0/$exit
      -- CP-element group 304: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_Sample/word_access_start/$exit
      -- CP-element group 304: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_Sample/$exit
      -- 
    ra_3215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1234_load_0_ack_0, ack => testConfigure_CP_0_elements(304)); -- 
    -- CP-element group 305:  transition  input  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	401 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (12) 
      -- CP-element group 305: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1238_Sample/rr
      -- CP-element group 305: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1238_Sample/$entry
      -- CP-element group 305: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_update_completed_
      -- CP-element group 305: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1238_sample_start_
      -- CP-element group 305: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_Update/ptr_deref_1234_Merge/merge_ack
      -- CP-element group 305: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_Update/ptr_deref_1234_Merge/merge_req
      -- CP-element group 305: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_Update/ptr_deref_1234_Merge/$exit
      -- CP-element group 305: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_Update/ptr_deref_1234_Merge/$entry
      -- CP-element group 305: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_Update/word_access_complete/word_0/ca
      -- CP-element group 305: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_Update/word_access_complete/word_0/$exit
      -- CP-element group 305: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_Update/word_access_complete/$exit
      -- CP-element group 305: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_Update/$exit
      -- 
    ca_3226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1234_load_0_ack_1, ack => testConfigure_CP_0_elements(305)); -- 
    rr_3239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(305), ack => type_cast_1238_inst_req_0); -- 
    -- CP-element group 306:  transition  input  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1238_Sample/ra
      -- CP-element group 306: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1238_Sample/$exit
      -- CP-element group 306: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1238_sample_completed_
      -- 
    ra_3240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_0, ack => testConfigure_CP_0_elements(306)); -- 
    -- CP-element group 307:  transition  input  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	401 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	312 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1238_Update/ca
      -- CP-element group 307: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1238_Update/$exit
      -- CP-element group 307: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1238_update_completed_
      -- 
    ca_3245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_1, ack => testConfigure_CP_0_elements(307)); -- 
    -- CP-element group 308:  transition  input  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	401 
    -- CP-element group 308: successors 
    -- CP-element group 308:  members (5) 
      -- CP-element group 308: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_sample_completed_
      -- CP-element group 308: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_Sample/word_access_start/word_0/ra
      -- CP-element group 308: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_Sample/word_access_start/word_0/$exit
      -- CP-element group 308: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_Sample/word_access_start/$exit
      -- CP-element group 308: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_Sample/$exit
      -- 
    ra_3279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1250_load_0_ack_0, ack => testConfigure_CP_0_elements(308)); -- 
    -- CP-element group 309:  transition  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	401 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (12) 
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_update_completed_
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_Update/word_access_complete/word_0/$exit
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_Update/word_access_complete/$exit
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_Update/$exit
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1254_Sample/rr
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1254_Sample/$entry
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1254_sample_start_
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_Update/ptr_deref_1250_Merge/merge_ack
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_Update/ptr_deref_1250_Merge/merge_req
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_Update/ptr_deref_1250_Merge/$exit
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_Update/ptr_deref_1250_Merge/$entry
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_Update/word_access_complete/word_0/ca
      -- 
    ca_3290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1250_load_0_ack_1, ack => testConfigure_CP_0_elements(309)); -- 
    rr_3303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(309), ack => type_cast_1254_inst_req_0); -- 
    -- CP-element group 310:  transition  input  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1254_Sample/ra
      -- CP-element group 310: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1254_Sample/$exit
      -- CP-element group 310: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1254_sample_completed_
      -- 
    ra_3304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1254_inst_ack_0, ack => testConfigure_CP_0_elements(310)); -- 
    -- CP-element group 311:  transition  input  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	401 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1254_Update/ca
      -- CP-element group 311: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1254_Update/$exit
      -- CP-element group 311: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1254_update_completed_
      -- 
    ca_3309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1254_inst_ack_1, ack => testConfigure_CP_0_elements(311)); -- 
    -- CP-element group 312:  branch  join  transition  place  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	303 
    -- CP-element group 312: 	307 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312: 	314 
    -- CP-element group 312:  members (10) 
      -- CP-element group 312: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271__exit__
      -- CP-element group 312: 	 branch_block_stmt_34/if_stmt_1272__entry__
      -- CP-element group 312: 	 branch_block_stmt_34/R_cmp281292_1273_place
      -- CP-element group 312: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/$exit
      -- CP-element group 312: 	 branch_block_stmt_34/if_stmt_1272_else_link/$entry
      -- CP-element group 312: 	 branch_block_stmt_34/if_stmt_1272_if_link/$entry
      -- CP-element group 312: 	 branch_block_stmt_34/if_stmt_1272_eval_test/branch_req
      -- CP-element group 312: 	 branch_block_stmt_34/if_stmt_1272_eval_test/$exit
      -- CP-element group 312: 	 branch_block_stmt_34/if_stmt_1272_eval_test/$entry
      -- CP-element group 312: 	 branch_block_stmt_34/if_stmt_1272_dead_link/$entry
      -- 
    branch_req_3317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(312), ack => if_stmt_1272_branch_req_0); -- 
    testConfigure_cp_element_group_312: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_312"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(303) & testConfigure_CP_0_elements(307) & testConfigure_CP_0_elements(311);
      gj_testConfigure_cp_element_group_312 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(312), clk => clk, reset => reset); --
    end block;
    -- CP-element group 313:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	315 
    -- CP-element group 313: 	316 
    -- CP-element group 313:  members (18) 
      -- CP-element group 313: 	 branch_block_stmt_34/merge_stmt_1278__exit__
      -- CP-element group 313: 	 branch_block_stmt_34/assign_stmt_1284_to_assign_stmt_1313__entry__
      -- CP-element group 313: 	 branch_block_stmt_34/forx_xend267_bbx_xnph
      -- CP-element group 313: 	 branch_block_stmt_34/assign_stmt_1284_to_assign_stmt_1313/type_cast_1299_Update/cr
      -- CP-element group 313: 	 branch_block_stmt_34/assign_stmt_1284_to_assign_stmt_1313/type_cast_1299_Update/$entry
      -- CP-element group 313: 	 branch_block_stmt_34/assign_stmt_1284_to_assign_stmt_1313/type_cast_1299_Sample/rr
      -- CP-element group 313: 	 branch_block_stmt_34/assign_stmt_1284_to_assign_stmt_1313/type_cast_1299_Sample/$entry
      -- CP-element group 313: 	 branch_block_stmt_34/assign_stmt_1284_to_assign_stmt_1313/type_cast_1299_update_start_
      -- CP-element group 313: 	 branch_block_stmt_34/assign_stmt_1284_to_assign_stmt_1313/type_cast_1299_sample_start_
      -- CP-element group 313: 	 branch_block_stmt_34/assign_stmt_1284_to_assign_stmt_1313/$entry
      -- CP-element group 313: 	 branch_block_stmt_34/if_stmt_1272_if_link/if_choice_transition
      -- CP-element group 313: 	 branch_block_stmt_34/if_stmt_1272_if_link/$exit
      -- CP-element group 313: 	 branch_block_stmt_34/forx_xend267_bbx_xnph_PhiReq/$entry
      -- CP-element group 313: 	 branch_block_stmt_34/forx_xend267_bbx_xnph_PhiReq/$exit
      -- CP-element group 313: 	 branch_block_stmt_34/merge_stmt_1278_PhiReqMerge
      -- CP-element group 313: 	 branch_block_stmt_34/merge_stmt_1278_PhiAck/$entry
      -- CP-element group 313: 	 branch_block_stmt_34/merge_stmt_1278_PhiAck/$exit
      -- CP-element group 313: 	 branch_block_stmt_34/merge_stmt_1278_PhiAck/dummy
      -- 
    if_choice_transition_3322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1272_branch_ack_1, ack => testConfigure_CP_0_elements(313)); -- 
    cr_3344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(313), ack => type_cast_1299_inst_req_1); -- 
    rr_3339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(313), ack => type_cast_1299_inst_req_0); -- 
    -- CP-element group 314:  transition  place  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	312 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	408 
    -- CP-element group 314:  members (5) 
      -- CP-element group 314: 	 branch_block_stmt_34/forx_xend267_forx_xend290
      -- CP-element group 314: 	 branch_block_stmt_34/if_stmt_1272_else_link/else_choice_transition
      -- CP-element group 314: 	 branch_block_stmt_34/if_stmt_1272_else_link/$exit
      -- CP-element group 314: 	 branch_block_stmt_34/forx_xend267_forx_xend290_PhiReq/$entry
      -- CP-element group 314: 	 branch_block_stmt_34/forx_xend267_forx_xend290_PhiReq/$exit
      -- 
    else_choice_transition_3326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1272_branch_ack_0, ack => testConfigure_CP_0_elements(314)); -- 
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	313 
    -- CP-element group 315: successors 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_34/assign_stmt_1284_to_assign_stmt_1313/type_cast_1299_Sample/ra
      -- CP-element group 315: 	 branch_block_stmt_34/assign_stmt_1284_to_assign_stmt_1313/type_cast_1299_Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_34/assign_stmt_1284_to_assign_stmt_1313/type_cast_1299_sample_completed_
      -- 
    ra_3340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1299_inst_ack_0, ack => testConfigure_CP_0_elements(315)); -- 
    -- CP-element group 316:  transition  place  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	313 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	402 
    -- CP-element group 316:  members (9) 
      -- CP-element group 316: 	 branch_block_stmt_34/assign_stmt_1284_to_assign_stmt_1313__exit__
      -- CP-element group 316: 	 branch_block_stmt_34/bbx_xnph_forx_xbody283
      -- CP-element group 316: 	 branch_block_stmt_34/assign_stmt_1284_to_assign_stmt_1313/type_cast_1299_Update/ca
      -- CP-element group 316: 	 branch_block_stmt_34/assign_stmt_1284_to_assign_stmt_1313/type_cast_1299_Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_34/assign_stmt_1284_to_assign_stmt_1313/type_cast_1299_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_34/assign_stmt_1284_to_assign_stmt_1313/$exit
      -- CP-element group 316: 	 branch_block_stmt_34/bbx_xnph_forx_xbody283_PhiReq/$entry
      -- CP-element group 316: 	 branch_block_stmt_34/bbx_xnph_forx_xbody283_PhiReq/phi_stmt_1316/$entry
      -- CP-element group 316: 	 branch_block_stmt_34/bbx_xnph_forx_xbody283_PhiReq/phi_stmt_1316/phi_stmt_1316_sources/$entry
      -- 
    ca_3345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1299_inst_ack_1, ack => testConfigure_CP_0_elements(316)); -- 
    -- CP-element group 317:  transition  input  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	407 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	323 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_final_index_sum_regn_sample_complete
      -- CP-element group 317: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_final_index_sum_regn_Sample/$exit
      -- CP-element group 317: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_final_index_sum_regn_Sample/ack
      -- 
    ack_3374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1328_index_offset_ack_0, ack => testConfigure_CP_0_elements(317)); -- 
    -- CP-element group 318:  transition  input  output  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	407 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (11) 
      -- CP-element group 318: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/addr_of_1329_request/$entry
      -- CP-element group 318: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_final_index_sum_regn_Update/$exit
      -- CP-element group 318: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_final_index_sum_regn_Update/ack
      -- CP-element group 318: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_base_plus_offset/$entry
      -- CP-element group 318: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_base_plus_offset/$exit
      -- CP-element group 318: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_base_plus_offset/sum_rename_req
      -- CP-element group 318: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_base_plus_offset/sum_rename_ack
      -- CP-element group 318: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_offset_calculated
      -- CP-element group 318: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_root_address_calculated
      -- CP-element group 318: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/addr_of_1329_sample_start_
      -- CP-element group 318: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/addr_of_1329_request/req
      -- 
    ack_3379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1328_index_offset_ack_1, ack => testConfigure_CP_0_elements(318)); -- 
    req_3388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(318), ack => addr_of_1329_final_reg_req_0); -- 
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/addr_of_1329_request/$exit
      -- CP-element group 319: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/addr_of_1329_sample_completed_
      -- CP-element group 319: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/addr_of_1329_request/ack
      -- 
    ack_3389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1329_final_reg_ack_0, ack => testConfigure_CP_0_elements(319)); -- 
    -- CP-element group 320:  join  fork  transition  input  output  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	407 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	321 
    -- CP-element group 320:  members (28) 
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_Sample/word_access_start/word_0/rr
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/addr_of_1329_update_completed_
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_Sample/word_access_start/word_0/$entry
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_Sample/word_access_start/$entry
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_Sample/ptr_deref_1332_Split/split_ack
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_Sample/ptr_deref_1332_Split/split_req
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_Sample/ptr_deref_1332_Split/$exit
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_Sample/ptr_deref_1332_Split/$entry
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_Sample/$entry
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_word_addrgen/root_register_ack
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_word_addrgen/root_register_req
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_word_addrgen/$exit
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_word_addrgen/$entry
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_base_plus_offset/sum_rename_ack
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_base_plus_offset/sum_rename_req
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_base_plus_offset/$exit
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_base_plus_offset/$entry
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_base_addr_resize/base_resize_ack
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_base_addr_resize/base_resize_req
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_base_addr_resize/$exit
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_base_addr_resize/$entry
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_base_address_resized
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_root_address_calculated
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_word_address_calculated
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_base_address_calculated
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_sample_start_
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/addr_of_1329_complete/ack
      -- CP-element group 320: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/addr_of_1329_complete/$exit
      -- 
    ack_3394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1329_final_reg_ack_1, ack => testConfigure_CP_0_elements(320)); -- 
    rr_3432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(320), ack => ptr_deref_1332_store_0_req_0); -- 
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	320 
    -- CP-element group 321: successors 
    -- CP-element group 321:  members (5) 
      -- CP-element group 321: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_Sample/word_access_start/word_0/ra
      -- CP-element group 321: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_Sample/word_access_start/word_0/$exit
      -- CP-element group 321: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_Sample/word_access_start/$exit
      -- CP-element group 321: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_Sample/$exit
      -- CP-element group 321: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_sample_completed_
      -- 
    ra_3433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1332_store_0_ack_0, ack => testConfigure_CP_0_elements(321)); -- 
    -- CP-element group 322:  transition  input  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	407 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (5) 
      -- CP-element group 322: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_Update/word_access_complete/word_0/$exit
      -- CP-element group 322: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_Update/word_access_complete/word_0/ca
      -- CP-element group 322: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_Update/word_access_complete/$exit
      -- CP-element group 322: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_Update/$exit
      -- CP-element group 322: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_update_completed_
      -- 
    ca_3444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1332_store_0_ack_1, ack => testConfigure_CP_0_elements(322)); -- 
    -- CP-element group 323:  branch  join  transition  place  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	317 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323: 	325 
    -- CP-element group 323:  members (10) 
      -- CP-element group 323: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346__exit__
      -- CP-element group 323: 	 branch_block_stmt_34/if_stmt_1347__entry__
      -- CP-element group 323: 	 branch_block_stmt_34/R_exitcond5_1348_place
      -- CP-element group 323: 	 branch_block_stmt_34/if_stmt_1347_dead_link/$entry
      -- CP-element group 323: 	 branch_block_stmt_34/if_stmt_1347_eval_test/$entry
      -- CP-element group 323: 	 branch_block_stmt_34/if_stmt_1347_eval_test/$exit
      -- CP-element group 323: 	 branch_block_stmt_34/if_stmt_1347_eval_test/branch_req
      -- CP-element group 323: 	 branch_block_stmt_34/if_stmt_1347_if_link/$entry
      -- CP-element group 323: 	 branch_block_stmt_34/if_stmt_1347_else_link/$entry
      -- CP-element group 323: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/$exit
      -- 
    branch_req_3452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(323), ack => if_stmt_1347_branch_req_0); -- 
    testConfigure_cp_element_group_323: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_323"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(317) & testConfigure_CP_0_elements(322);
      gj_testConfigure_cp_element_group_323 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(323), clk => clk, reset => reset); --
    end block;
    -- CP-element group 324:  merge  transition  place  input  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	408 
    -- CP-element group 324:  members (13) 
      -- CP-element group 324: 	 branch_block_stmt_34/merge_stmt_1353__exit__
      -- CP-element group 324: 	 branch_block_stmt_34/forx_xend290x_xloopexit_forx_xend290
      -- CP-element group 324: 	 branch_block_stmt_34/forx_xbody283_forx_xend290x_xloopexit
      -- CP-element group 324: 	 branch_block_stmt_34/if_stmt_1347_if_link/$exit
      -- CP-element group 324: 	 branch_block_stmt_34/if_stmt_1347_if_link/if_choice_transition
      -- CP-element group 324: 	 branch_block_stmt_34/forx_xbody283_forx_xend290x_xloopexit_PhiReq/$entry
      -- CP-element group 324: 	 branch_block_stmt_34/forx_xbody283_forx_xend290x_xloopexit_PhiReq/$exit
      -- CP-element group 324: 	 branch_block_stmt_34/merge_stmt_1353_PhiReqMerge
      -- CP-element group 324: 	 branch_block_stmt_34/merge_stmt_1353_PhiAck/$entry
      -- CP-element group 324: 	 branch_block_stmt_34/merge_stmt_1353_PhiAck/$exit
      -- CP-element group 324: 	 branch_block_stmt_34/merge_stmt_1353_PhiAck/dummy
      -- CP-element group 324: 	 branch_block_stmt_34/forx_xend290x_xloopexit_forx_xend290_PhiReq/$entry
      -- CP-element group 324: 	 branch_block_stmt_34/forx_xend290x_xloopexit_forx_xend290_PhiReq/$exit
      -- 
    if_choice_transition_3457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1347_branch_ack_1, ack => testConfigure_CP_0_elements(324)); -- 
    -- CP-element group 325:  fork  transition  place  input  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	323 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	403 
    -- CP-element group 325: 	404 
    -- CP-element group 325:  members (12) 
      -- CP-element group 325: 	 branch_block_stmt_34/forx_xbody283_forx_xbody283
      -- CP-element group 325: 	 branch_block_stmt_34/if_stmt_1347_else_link/$exit
      -- CP-element group 325: 	 branch_block_stmt_34/if_stmt_1347_else_link/else_choice_transition
      -- CP-element group 325: 	 branch_block_stmt_34/forx_xbody283_forx_xbody283_PhiReq/$entry
      -- CP-element group 325: 	 branch_block_stmt_34/forx_xbody283_forx_xbody283_PhiReq/phi_stmt_1316/$entry
      -- CP-element group 325: 	 branch_block_stmt_34/forx_xbody283_forx_xbody283_PhiReq/phi_stmt_1316/phi_stmt_1316_sources/$entry
      -- CP-element group 325: 	 branch_block_stmt_34/forx_xbody283_forx_xbody283_PhiReq/phi_stmt_1316/phi_stmt_1316_sources/type_cast_1322/$entry
      -- CP-element group 325: 	 branch_block_stmt_34/forx_xbody283_forx_xbody283_PhiReq/phi_stmt_1316/phi_stmt_1316_sources/type_cast_1322/SplitProtocol/$entry
      -- CP-element group 325: 	 branch_block_stmt_34/forx_xbody283_forx_xbody283_PhiReq/phi_stmt_1316/phi_stmt_1316_sources/type_cast_1322/SplitProtocol/Sample/$entry
      -- CP-element group 325: 	 branch_block_stmt_34/forx_xbody283_forx_xbody283_PhiReq/phi_stmt_1316/phi_stmt_1316_sources/type_cast_1322/SplitProtocol/Sample/rr
      -- CP-element group 325: 	 branch_block_stmt_34/forx_xbody283_forx_xbody283_PhiReq/phi_stmt_1316/phi_stmt_1316_sources/type_cast_1322/SplitProtocol/Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_34/forx_xbody283_forx_xbody283_PhiReq/phi_stmt_1316/phi_stmt_1316_sources/type_cast_1322/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1347_branch_ack_0, ack => testConfigure_CP_0_elements(325)); -- 
    rr_4080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(325), ack => type_cast_1322_inst_req_0); -- 
    cr_4085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(325), ack => type_cast_1322_inst_req_1); -- 
    -- CP-element group 326:  transition  input  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	51 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	328 
    -- CP-element group 326:  members (2) 
      -- CP-element group 326: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_103/phi_stmt_103_sources/type_cast_106/SplitProtocol/Sample/ra
      -- CP-element group 326: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_103/phi_stmt_103_sources/type_cast_106/SplitProtocol/Sample/$exit
      -- 
    ra_3498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_106_inst_ack_0, ack => testConfigure_CP_0_elements(326)); -- 
    -- CP-element group 327:  transition  input  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	51 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (2) 
      -- CP-element group 327: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_103/phi_stmt_103_sources/type_cast_106/SplitProtocol/Update/ca
      -- CP-element group 327: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_103/phi_stmt_103_sources/type_cast_106/SplitProtocol/Update/$exit
      -- 
    ca_3503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_106_inst_ack_1, ack => testConfigure_CP_0_elements(327)); -- 
    -- CP-element group 328:  join  transition  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	326 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	332 
    -- CP-element group 328:  members (5) 
      -- CP-element group 328: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_103/phi_stmt_103_req
      -- CP-element group 328: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_103/phi_stmt_103_sources/type_cast_106/SplitProtocol/$exit
      -- CP-element group 328: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_103/phi_stmt_103_sources/type_cast_106/$exit
      -- CP-element group 328: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_103/phi_stmt_103_sources/$exit
      -- CP-element group 328: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_103/$exit
      -- 
    phi_stmt_103_req_3504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_103_req_3504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(328), ack => phi_stmt_103_req_0); -- 
    testConfigure_cp_element_group_328: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_328"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(326) & testConfigure_CP_0_elements(327);
      gj_testConfigure_cp_element_group_328 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(328), clk => clk, reset => reset); --
    end block;
    -- CP-element group 329:  transition  input  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	51 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	331 
    -- CP-element group 329:  members (2) 
      -- CP-element group 329: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_115/SplitProtocol/Sample/$exit
      -- CP-element group 329: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_115/SplitProtocol/Sample/ra
      -- 
    ra_3521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_115_inst_ack_0, ack => testConfigure_CP_0_elements(329)); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	51 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	331 
    -- CP-element group 330:  members (2) 
      -- CP-element group 330: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_115/SplitProtocol/Update/$exit
      -- CP-element group 330: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_115/SplitProtocol/Update/ca
      -- 
    ca_3526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_115_inst_ack_1, ack => testConfigure_CP_0_elements(330)); -- 
    -- CP-element group 331:  join  transition  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	329 
    -- CP-element group 331: 	330 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (5) 
      -- CP-element group 331: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_115/SplitProtocol/$exit
      -- CP-element group 331: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_115/$exit
      -- CP-element group 331: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/$exit
      -- CP-element group 331: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_110/$exit
      -- CP-element group 331: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_req
      -- 
    phi_stmt_110_req_3527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_110_req_3527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(331), ack => phi_stmt_110_req_1); -- 
    testConfigure_cp_element_group_331: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_331"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(329) & testConfigure_CP_0_elements(330);
      gj_testConfigure_cp_element_group_331 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(331), clk => clk, reset => reset); --
    end block;
    -- CP-element group 332:  join  transition  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	328 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	338 
    -- CP-element group 332:  members (1) 
      -- CP-element group 332: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_332: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_332"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(328) & testConfigure_CP_0_elements(331);
      gj_testConfigure_cp_element_group_332 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(332), clk => clk, reset => reset); --
    end block;
    -- CP-element group 333:  transition  output  delay-element  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	23 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	337 
    -- CP-element group 333:  members (4) 
      -- CP-element group 333: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_103/phi_stmt_103_req
      -- CP-element group 333: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_103/phi_stmt_103_sources/type_cast_109_konst_delay_trans
      -- CP-element group 333: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_103/phi_stmt_103_sources/$exit
      -- CP-element group 333: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_103/$exit
      -- 
    phi_stmt_103_req_3538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_103_req_3538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(333), ack => phi_stmt_103_req_1); -- 
    -- Element group testConfigure_CP_0_elements(333) is a control-delay.
    cp_element_333_delay: control_delay_element  generic map(name => " 333_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(23), ack => testConfigure_CP_0_elements(333), clk => clk, reset =>reset);
    -- CP-element group 334:  transition  input  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	23 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	336 
    -- CP-element group 334:  members (2) 
      -- CP-element group 334: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_113/SplitProtocol/Sample/ra
      -- CP-element group 334: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_113/SplitProtocol/Sample/$exit
      -- 
    ra_3555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_113_inst_ack_0, ack => testConfigure_CP_0_elements(334)); -- 
    -- CP-element group 335:  transition  input  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	23 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (2) 
      -- CP-element group 335: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_113/SplitProtocol/Update/ca
      -- CP-element group 335: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_113/SplitProtocol/Update/$exit
      -- 
    ca_3560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_113_inst_ack_1, ack => testConfigure_CP_0_elements(335)); -- 
    -- CP-element group 336:  join  transition  output  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	334 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336:  members (5) 
      -- CP-element group 336: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_req
      -- CP-element group 336: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_113/SplitProtocol/$exit
      -- CP-element group 336: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/type_cast_113/$exit
      -- CP-element group 336: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_110/phi_stmt_110_sources/$exit
      -- CP-element group 336: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_110/$exit
      -- 
    phi_stmt_110_req_3561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_110_req_3561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(336), ack => phi_stmt_110_req_0); -- 
    testConfigure_cp_element_group_336: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_336"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(334) & testConfigure_CP_0_elements(335);
      gj_testConfigure_cp_element_group_336 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(336), clk => clk, reset => reset); --
    end block;
    -- CP-element group 337:  join  transition  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	333 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (1) 
      -- CP-element group 337: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_337: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_337"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(333) & testConfigure_CP_0_elements(336);
      gj_testConfigure_cp_element_group_337 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(337), clk => clk, reset => reset); --
    end block;
    -- CP-element group 338:  merge  fork  transition  place  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	332 
    -- CP-element group 338: 	337 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338: 	340 
    -- CP-element group 338:  members (2) 
      -- CP-element group 338: 	 branch_block_stmt_34/merge_stmt_102_PhiAck/$entry
      -- CP-element group 338: 	 branch_block_stmt_34/merge_stmt_102_PhiReqMerge
      -- 
    testConfigure_CP_0_elements(338) <= OrReduce(testConfigure_CP_0_elements(332) & testConfigure_CP_0_elements(337));
    -- CP-element group 339:  transition  input  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	338 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	341 
    -- CP-element group 339:  members (1) 
      -- CP-element group 339: 	 branch_block_stmt_34/merge_stmt_102_PhiAck/phi_stmt_103_ack
      -- 
    phi_stmt_103_ack_3566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_103_ack_0, ack => testConfigure_CP_0_elements(339)); -- 
    -- CP-element group 340:  transition  input  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	338 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (1) 
      -- CP-element group 340: 	 branch_block_stmt_34/merge_stmt_102_PhiAck/phi_stmt_110_ack
      -- 
    phi_stmt_110_ack_3567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_110_ack_0, ack => testConfigure_CP_0_elements(340)); -- 
    -- CP-element group 341:  join  fork  transition  place  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	339 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	41 
    -- CP-element group 341: 	43 
    -- CP-element group 341: 	24 
    -- CP-element group 341: 	25 
    -- CP-element group 341: 	26 
    -- CP-element group 341: 	27 
    -- CP-element group 341: 	29 
    -- CP-element group 341: 	31 
    -- CP-element group 341: 	32 
    -- CP-element group 341: 	35 
    -- CP-element group 341: 	38 
    -- CP-element group 341: 	39 
    -- CP-element group 341: 	47 
    -- CP-element group 341:  members (72) 
      -- CP-element group 341: 	 branch_block_stmt_34/merge_stmt_102__exit__
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194__entry__
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/addr_of_132_update_start_
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_index_resized_1
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_index_scaled_1
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_index_computed_1
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_index_resize_1/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_index_resize_1/$exit
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_index_resize_1/index_resize_req
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_index_resize_1/index_resize_ack
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_index_scale_1/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_index_scale_1/$exit
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_index_scale_1/scale_rename_req
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_125_sample_start_
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_125_update_start_
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_125_Sample/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_125_Sample/rr
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_125_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_125_Update/cr
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_index_scale_1/scale_rename_ack
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_final_index_sum_regn_update_start
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_final_index_sum_regn_Sample/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_final_index_sum_regn_Sample/req
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_final_index_sum_regn_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/array_obj_ref_131_final_index_sum_regn_Update/req
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/addr_of_132_complete/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/addr_of_132_complete/req
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_update_start_
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_Update/word_access_complete/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_Update/word_access_complete/word_0/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_135_Update/word_access_complete/word_0/cr
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_145_sample_start_
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_145_Sample/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/RPIPE_ConvTranspose_input_pipe_145_Sample/rr
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_149_update_start_
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_149_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_149_Update/cr
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_update_start_
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_Update/word_access_complete/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_Update/word_access_complete/word_0/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_157_Update/word_access_complete/word_0/cr
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_update_start_
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_base_address_calculated
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_word_address_calculated
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_root_address_calculated
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_base_address_resized
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_base_addr_resize/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_base_addr_resize/$exit
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_base_addr_resize/base_resize_req
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_base_addr_resize/base_resize_ack
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_base_plus_offset/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_base_plus_offset/$exit
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_base_plus_offset/sum_rename_req
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_base_plus_offset/sum_rename_ack
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_word_addrgen/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_word_addrgen/$exit
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_word_addrgen/root_register_req
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_word_addrgen/root_register_ack
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_Update/word_access_complete/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_Update/word_access_complete/word_0/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/ptr_deref_174_Update/word_access_complete/word_0/cr
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_178_update_start_
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_178_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_178_Update/cr
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_193_update_start_
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_193_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_34/assign_stmt_122_to_assign_stmt_194/type_cast_193_Update/cr
      -- CP-element group 341: 	 branch_block_stmt_34/merge_stmt_102_PhiAck/$exit
      -- 
    rr_325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(341), ack => type_cast_125_inst_req_0); -- 
    cr_330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(341), ack => type_cast_125_inst_req_1); -- 
    req_356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(341), ack => array_obj_ref_131_index_offset_req_0); -- 
    req_361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(341), ack => array_obj_ref_131_index_offset_req_1); -- 
    req_376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(341), ack => addr_of_132_final_reg_req_1); -- 
    cr_426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(341), ack => ptr_deref_135_store_0_req_1); -- 
    rr_435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(341), ack => RPIPE_ConvTranspose_input_pipe_145_inst_req_0); -- 
    cr_454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(341), ack => type_cast_149_inst_req_1); -- 
    cr_504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(341), ack => ptr_deref_157_store_0_req_1); -- 
    cr_549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(341), ack => ptr_deref_174_load_0_req_1); -- 
    cr_568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(341), ack => type_cast_178_inst_req_1); -- 
    cr_596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(341), ack => type_cast_193_inst_req_1); -- 
    testConfigure_cp_element_group_341: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_341"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(339) & testConfigure_CP_0_elements(340);
      gj_testConfigure_cp_element_group_341 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(341), clk => clk, reset => reset); --
    end block;
    -- CP-element group 342:  transition  input  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	52 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	344 
    -- CP-element group 342:  members (2) 
      -- CP-element group 342: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_202/phi_stmt_202_sources/type_cast_205/SplitProtocol/Sample/$exit
      -- CP-element group 342: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_202/phi_stmt_202_sources/type_cast_205/SplitProtocol/Sample/ra
      -- 
    ra_3591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_205_inst_ack_0, ack => testConfigure_CP_0_elements(342)); -- 
    -- CP-element group 343:  transition  input  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	52 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343:  members (2) 
      -- CP-element group 343: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_202/phi_stmt_202_sources/type_cast_205/SplitProtocol/Update/$exit
      -- CP-element group 343: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_202/phi_stmt_202_sources/type_cast_205/SplitProtocol/Update/ca
      -- 
    ca_3596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_205_inst_ack_1, ack => testConfigure_CP_0_elements(343)); -- 
    -- CP-element group 344:  join  transition  place  output  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	342 
    -- CP-element group 344: 	343 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	345 
    -- CP-element group 344:  members (8) 
      -- CP-element group 344: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_202/phi_stmt_202_sources/type_cast_205/SplitProtocol/$exit
      -- CP-element group 344: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_202/phi_stmt_202_sources/type_cast_205/$exit
      -- CP-element group 344: 	 branch_block_stmt_34/merge_stmt_201_PhiAck/$entry
      -- CP-element group 344: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_202/phi_stmt_202_sources/$exit
      -- CP-element group 344: 	 branch_block_stmt_34/merge_stmt_201_PhiReqMerge
      -- CP-element group 344: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_202/$exit
      -- CP-element group 344: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 344: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_202/phi_stmt_202_req
      -- 
    phi_stmt_202_req_3597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_202_req_3597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(344), ack => phi_stmt_202_req_0); -- 
    testConfigure_cp_element_group_344: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_344"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(342) & testConfigure_CP_0_elements(343);
      gj_testConfigure_cp_element_group_344 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(344), clk => clk, reset => reset); --
    end block;
    -- CP-element group 345:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	344 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	349 
    -- CP-element group 345: 	350 
    -- CP-element group 345:  members (13) 
      -- CP-element group 345: 	 branch_block_stmt_34/merge_stmt_201__exit__
      -- CP-element group 345: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend
      -- CP-element group 345: 	 branch_block_stmt_34/merge_stmt_201_PhiAck/$exit
      -- CP-element group 345: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/$entry
      -- CP-element group 345: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_209/$entry
      -- CP-element group 345: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 345: 	 branch_block_stmt_34/merge_stmt_201_PhiAck/phi_stmt_202_ack
      -- CP-element group 345: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_214/$entry
      -- CP-element group 345: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_214/SplitProtocol/$entry
      -- CP-element group 345: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_214/SplitProtocol/Sample/$entry
      -- CP-element group 345: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_214/SplitProtocol/Sample/rr
      -- CP-element group 345: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_214/SplitProtocol/Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_214/SplitProtocol/Update/cr
      -- 
    phi_stmt_202_ack_3602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_202_ack_0, ack => testConfigure_CP_0_elements(345)); -- 
    rr_3647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(345), ack => type_cast_214_inst_req_0); -- 
    cr_3652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(345), ack => type_cast_214_inst_req_1); -- 
    -- CP-element group 346:  transition  input  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	22 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	348 
    -- CP-element group 346:  members (2) 
      -- CP-element group 346: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_212/SplitProtocol/Sample/ra
      -- CP-element group 346: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_212/SplitProtocol/Sample/$exit
      -- 
    ra_3622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_212_inst_ack_0, ack => testConfigure_CP_0_elements(346)); -- 
    -- CP-element group 347:  transition  input  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	22 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (2) 
      -- CP-element group 347: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_212/SplitProtocol/Update/$exit
      -- CP-element group 347: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_212/SplitProtocol/Update/ca
      -- 
    ca_3627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_212_inst_ack_1, ack => testConfigure_CP_0_elements(347)); -- 
    -- CP-element group 348:  join  transition  output  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	346 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	352 
    -- CP-element group 348:  members (6) 
      -- CP-element group 348: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/$exit
      -- CP-element group 348: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_209/$exit
      -- CP-element group 348: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_req
      -- CP-element group 348: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/$exit
      -- CP-element group 348: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_212/SplitProtocol/$exit
      -- CP-element group 348: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_212/$exit
      -- 
    phi_stmt_209_req_3628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_209_req_3628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(348), ack => phi_stmt_209_req_0); -- 
    testConfigure_cp_element_group_348: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_348"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(346) & testConfigure_CP_0_elements(347);
      gj_testConfigure_cp_element_group_348 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(348), clk => clk, reset => reset); --
    end block;
    -- CP-element group 349:  transition  input  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	345 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	351 
    -- CP-element group 349:  members (2) 
      -- CP-element group 349: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_214/SplitProtocol/Sample/$exit
      -- CP-element group 349: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_214/SplitProtocol/Sample/ra
      -- 
    ra_3648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_214_inst_ack_0, ack => testConfigure_CP_0_elements(349)); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	345 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	351 
    -- CP-element group 350:  members (2) 
      -- CP-element group 350: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_214/SplitProtocol/Update/$exit
      -- CP-element group 350: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_214/SplitProtocol/Update/ca
      -- 
    ca_3653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_214_inst_ack_1, ack => testConfigure_CP_0_elements(350)); -- 
    -- CP-element group 351:  join  transition  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	349 
    -- CP-element group 351: 	350 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (6) 
      -- CP-element group 351: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_209/$exit
      -- CP-element group 351: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- CP-element group 351: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/$exit
      -- CP-element group 351: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_214/$exit
      -- CP-element group 351: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_sources/type_cast_214/SplitProtocol/$exit
      -- CP-element group 351: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_209/phi_stmt_209_req
      -- 
    phi_stmt_209_req_3654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_209_req_3654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(351), ack => phi_stmt_209_req_1); -- 
    testConfigure_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(349) & testConfigure_CP_0_elements(350);
      gj_testConfigure_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  merge  transition  place  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	348 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (2) 
      -- CP-element group 352: 	 branch_block_stmt_34/merge_stmt_208_PhiReqMerge
      -- CP-element group 352: 	 branch_block_stmt_34/merge_stmt_208_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(352) <= OrReduce(testConfigure_CP_0_elements(348) & testConfigure_CP_0_elements(351));
    -- CP-element group 353:  join  fork  transition  place  input  output  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	53 
    -- CP-element group 353: 	54 
    -- CP-element group 353: 	55 
    -- CP-element group 353: 	58 
    -- CP-element group 353: 	59 
    -- CP-element group 353: 	61 
    -- CP-element group 353:  members (62) 
      -- CP-element group 353: 	 branch_block_stmt_34/merge_stmt_208__exit__
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259__entry__
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/$entry
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_sample_start_
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_update_start_
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_base_address_calculated
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_word_address_calculated
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_root_address_calculated
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_base_address_resized
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_base_addr_resize/$entry
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_base_addr_resize/$exit
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_base_addr_resize/base_resize_req
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_base_addr_resize/base_resize_ack
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_base_plus_offset/$entry
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_base_plus_offset/$exit
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_base_plus_offset/sum_rename_req
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_base_plus_offset/sum_rename_ack
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_word_addrgen/$entry
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_word_addrgen/$exit
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_word_addrgen/root_register_req
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_word_addrgen/root_register_ack
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_Sample/$entry
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_Sample/ptr_deref_223_Split/$entry
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_Sample/ptr_deref_223_Split/$exit
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_Sample/ptr_deref_223_Split/split_req
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_Sample/ptr_deref_223_Split/split_ack
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_Sample/word_access_start/$entry
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_Sample/word_access_start/word_0/$entry
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_Sample/word_access_start/word_0/rr
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_Update/$entry
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_Update/word_access_complete/$entry
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_Update/word_access_complete/word_0/$entry
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_223_Update/word_access_complete/word_0/cr
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/RPIPE_ConvTranspose_input_pipe_233_sample_start_
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/RPIPE_ConvTranspose_input_pipe_233_Sample/$entry
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/RPIPE_ConvTranspose_input_pipe_233_Sample/rr
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/type_cast_237_update_start_
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/type_cast_237_Update/$entry
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/type_cast_237_Update/cr
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_update_start_
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_base_address_calculated
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_word_address_calculated
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_root_address_calculated
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_base_address_resized
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_base_addr_resize/$entry
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_base_addr_resize/$exit
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_base_addr_resize/base_resize_req
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_base_addr_resize/base_resize_ack
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_base_plus_offset/$entry
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_base_plus_offset/$exit
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_base_plus_offset/sum_rename_req
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_base_plus_offset/sum_rename_ack
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_word_addrgen/$entry
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_word_addrgen/$exit
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_word_addrgen/root_register_req
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_word_addrgen/root_register_ack
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_Update/$entry
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_Update/word_access_complete/$entry
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_Update/word_access_complete/word_0/$entry
      -- CP-element group 353: 	 branch_block_stmt_34/assign_stmt_221_to_assign_stmt_259/ptr_deref_251_Update/word_access_complete/word_0/cr
      -- CP-element group 353: 	 branch_block_stmt_34/merge_stmt_208_PhiAck/$exit
      -- CP-element group 353: 	 branch_block_stmt_34/merge_stmt_208_PhiAck/phi_stmt_209_ack
      -- 
    phi_stmt_209_ack_3659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_209_ack_0, ack => testConfigure_CP_0_elements(353)); -- 
    rr_659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(353), ack => ptr_deref_223_store_0_req_0); -- 
    cr_670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(353), ack => ptr_deref_223_store_0_req_1); -- 
    rr_679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(353), ack => RPIPE_ConvTranspose_input_pipe_233_inst_req_0); -- 
    cr_698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(353), ack => type_cast_237_inst_req_1); -- 
    cr_748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(353), ack => ptr_deref_251_store_0_req_1); -- 
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	94 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	356 
    -- CP-element group 354:  members (2) 
      -- CP-element group 354: 	 branch_block_stmt_34/forx_xbody42_forx_xbody42_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_272/SplitProtocol/Sample/$exit
      -- CP-element group 354: 	 branch_block_stmt_34/forx_xbody42_forx_xbody42_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_272/SplitProtocol/Sample/ra
      -- 
    ra_3691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_272_inst_ack_0, ack => testConfigure_CP_0_elements(354)); -- 
    -- CP-element group 355:  transition  input  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	94 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (2) 
      -- CP-element group 355: 	 branch_block_stmt_34/forx_xbody42_forx_xbody42_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_272/SplitProtocol/Update/$exit
      -- CP-element group 355: 	 branch_block_stmt_34/forx_xbody42_forx_xbody42_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_272/SplitProtocol/Update/ca
      -- 
    ca_3696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_272_inst_ack_1, ack => testConfigure_CP_0_elements(355)); -- 
    -- CP-element group 356:  join  transition  output  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	354 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	358 
    -- CP-element group 356:  members (6) 
      -- CP-element group 356: 	 branch_block_stmt_34/forx_xbody42_forx_xbody42_PhiReq/$exit
      -- CP-element group 356: 	 branch_block_stmt_34/forx_xbody42_forx_xbody42_PhiReq/phi_stmt_269/$exit
      -- CP-element group 356: 	 branch_block_stmt_34/forx_xbody42_forx_xbody42_PhiReq/phi_stmt_269/phi_stmt_269_sources/$exit
      -- CP-element group 356: 	 branch_block_stmt_34/forx_xbody42_forx_xbody42_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_272/$exit
      -- CP-element group 356: 	 branch_block_stmt_34/forx_xbody42_forx_xbody42_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_272/SplitProtocol/$exit
      -- CP-element group 356: 	 branch_block_stmt_34/forx_xbody42_forx_xbody42_PhiReq/phi_stmt_269/phi_stmt_269_req
      -- 
    phi_stmt_269_req_3697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_269_req_3697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(356), ack => phi_stmt_269_req_0); -- 
    testConfigure_cp_element_group_356: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_356"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(354) & testConfigure_CP_0_elements(355);
      gj_testConfigure_cp_element_group_356 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(356), clk => clk, reset => reset); --
    end block;
    -- CP-element group 357:  transition  output  delay-element  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	65 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (5) 
      -- CP-element group 357: 	 branch_block_stmt_34/forx_xbody42x_xpreheader_forx_xbody42_PhiReq/$exit
      -- CP-element group 357: 	 branch_block_stmt_34/forx_xbody42x_xpreheader_forx_xbody42_PhiReq/phi_stmt_269/$exit
      -- CP-element group 357: 	 branch_block_stmt_34/forx_xbody42x_xpreheader_forx_xbody42_PhiReq/phi_stmt_269/phi_stmt_269_sources/$exit
      -- CP-element group 357: 	 branch_block_stmt_34/forx_xbody42x_xpreheader_forx_xbody42_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_275_konst_delay_trans
      -- CP-element group 357: 	 branch_block_stmt_34/forx_xbody42x_xpreheader_forx_xbody42_PhiReq/phi_stmt_269/phi_stmt_269_req
      -- 
    phi_stmt_269_req_3708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_269_req_3708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(357), ack => phi_stmt_269_req_1); -- 
    -- Element group testConfigure_CP_0_elements(357) is a control-delay.
    cp_element_357_delay: control_delay_element  generic map(name => " 357_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(65), ack => testConfigure_CP_0_elements(357), clk => clk, reset =>reset);
    -- CP-element group 358:  merge  transition  place  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	356 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (2) 
      -- CP-element group 358: 	 branch_block_stmt_34/merge_stmt_268_PhiReqMerge
      -- CP-element group 358: 	 branch_block_stmt_34/merge_stmt_268_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(358) <= OrReduce(testConfigure_CP_0_elements(356) & testConfigure_CP_0_elements(357));
    -- CP-element group 359:  fork  transition  place  input  output  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	66 
    -- CP-element group 359: 	67 
    -- CP-element group 359: 	68 
    -- CP-element group 359: 	69 
    -- CP-element group 359: 	71 
    -- CP-element group 359: 	72 
    -- CP-element group 359: 	75 
    -- CP-element group 359: 	78 
    -- CP-element group 359: 	82 
    -- CP-element group 359: 	85 
    -- CP-element group 359: 	86 
    -- CP-element group 359: 	88 
    -- CP-element group 359: 	90 
    -- CP-element group 359:  members (73) 
      -- CP-element group 359: 	 branch_block_stmt_34/merge_stmt_268__exit__
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353__entry__
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_285_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_285_Update/cr
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/addr_of_292_update_start_
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_index_resized_1
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_index_scaled_1
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_index_computed_1
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_index_resize_1/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_index_resize_1/$exit
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_index_resize_1/index_resize_req
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_index_resize_1/index_resize_ack
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_index_scale_1/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_index_scale_1/$exit
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_index_scale_1/scale_rename_req
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_index_scale_1/scale_rename_ack
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_285_sample_start_
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_285_update_start_
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_285_Sample/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_285_Sample/rr
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_final_index_sum_regn_update_start
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_final_index_sum_regn_Sample/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_final_index_sum_regn_Sample/req
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_final_index_sum_regn_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/array_obj_ref_291_final_index_sum_regn_Update/req
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/addr_of_292_complete/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/addr_of_292_complete/req
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_295_sample_start_
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_295_Sample/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/RPIPE_ConvTranspose_input_pipe_295_Sample/rr
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_299_update_start_
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_299_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_299_Update/cr
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_update_start_
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_Update/word_access_complete/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_Update/word_access_complete/word_0/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_302_Update/word_access_complete/word_0/cr
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_316_update_start_
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_316_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_316_Update/cr
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_update_start_
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_Update/word_access_complete/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_Update/word_access_complete/word_0/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_324_Update/word_access_complete/word_0/cr
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_update_start_
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_base_address_calculated
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_word_address_calculated
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_root_address_calculated
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_base_address_resized
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_base_addr_resize/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_base_addr_resize/$exit
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_base_addr_resize/base_resize_req
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_base_addr_resize/base_resize_ack
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_base_plus_offset/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_base_plus_offset/$exit
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_base_plus_offset/sum_rename_req
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_base_plus_offset/sum_rename_ack
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_word_addrgen/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_word_addrgen/$exit
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_word_addrgen/root_register_req
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_word_addrgen/root_register_ack
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_Update/word_access_complete/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_Update/word_access_complete/word_0/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/ptr_deref_341_Update/word_access_complete/word_0/cr
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_345_update_start_
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_345_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_34/assign_stmt_282_to_assign_stmt_353/type_cast_345_Update/cr
      -- CP-element group 359: 	 branch_block_stmt_34/merge_stmt_268_PhiAck/$exit
      -- CP-element group 359: 	 branch_block_stmt_34/merge_stmt_268_PhiAck/phi_stmt_269_ack
      -- 
    phi_stmt_269_ack_3713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_269_ack_0, ack => testConfigure_CP_0_elements(359)); -- 
    cr_785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(359), ack => type_cast_285_inst_req_1); -- 
    rr_780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(359), ack => type_cast_285_inst_req_0); -- 
    req_811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(359), ack => array_obj_ref_291_index_offset_req_0); -- 
    req_816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(359), ack => array_obj_ref_291_index_offset_req_1); -- 
    req_831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(359), ack => addr_of_292_final_reg_req_1); -- 
    rr_840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(359), ack => RPIPE_ConvTranspose_input_pipe_295_inst_req_0); -- 
    cr_859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(359), ack => type_cast_299_inst_req_1); -- 
    cr_909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(359), ack => ptr_deref_302_store_0_req_1); -- 
    cr_937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(359), ack => type_cast_316_inst_req_1); -- 
    cr_987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(359), ack => ptr_deref_324_store_0_req_1); -- 
    cr_1032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(359), ack => ptr_deref_341_load_0_req_1); -- 
    cr_1051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(359), ack => type_cast_345_inst_req_1); -- 
    -- CP-element group 360:  merge  fork  transition  place  output  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	64 
    -- CP-element group 360: 	95 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	96 
    -- CP-element group 360: 	99 
    -- CP-element group 360:  members (13) 
      -- CP-element group 360: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/RPIPE_ConvTranspose_input_pipe_364_Sample/rr
      -- CP-element group 360: 	 branch_block_stmt_34/merge_stmt_362__exit__
      -- CP-element group 360: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369__entry__
      -- CP-element group 360: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/type_cast_368_Update/cr
      -- CP-element group 360: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/RPIPE_ConvTranspose_input_pipe_364_Sample/$entry
      -- CP-element group 360: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/type_cast_368_Update/$entry
      -- CP-element group 360: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/type_cast_368_update_start_
      -- CP-element group 360: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/RPIPE_ConvTranspose_input_pipe_364_sample_start_
      -- CP-element group 360: 	 branch_block_stmt_34/assign_stmt_365_to_assign_stmt_369/$entry
      -- CP-element group 360: 	 branch_block_stmt_34/merge_stmt_362_PhiReqMerge
      -- CP-element group 360: 	 branch_block_stmt_34/merge_stmt_362_PhiAck/$entry
      -- CP-element group 360: 	 branch_block_stmt_34/merge_stmt_362_PhiAck/$exit
      -- CP-element group 360: 	 branch_block_stmt_34/merge_stmt_362_PhiAck/dummy
      -- 
    rr_1084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(360), ack => RPIPE_ConvTranspose_input_pipe_364_inst_req_0); -- 
    cr_1103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(360), ack => type_cast_368_inst_req_1); -- 
    testConfigure_CP_0_elements(360) <= OrReduce(testConfigure_CP_0_elements(64) & testConfigure_CP_0_elements(95));
    -- CP-element group 361:  transition  output  delay-element  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	99 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	365 
    -- CP-element group 361:  members (4) 
      -- CP-element group 361: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_372/$exit
      -- CP-element group 361: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_372/phi_stmt_372_sources/$exit
      -- CP-element group 361: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_372/phi_stmt_372_sources/type_cast_376_konst_delay_trans
      -- CP-element group 361: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_372/phi_stmt_372_req
      -- 
    phi_stmt_372_req_3747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_372_req_3747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(361), ack => phi_stmt_372_req_0); -- 
    -- Element group testConfigure_CP_0_elements(361) is a control-delay.
    cp_element_361_delay: control_delay_element  generic map(name => " 361_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(99), ack => testConfigure_CP_0_elements(361), clk => clk, reset =>reset);
    -- CP-element group 362:  transition  input  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	99 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	364 
    -- CP-element group 362:  members (2) 
      -- CP-element group 362: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_382/SplitProtocol/Sample/$exit
      -- CP-element group 362: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_382/SplitProtocol/Sample/ra
      -- 
    ra_3764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_382_inst_ack_0, ack => testConfigure_CP_0_elements(362)); -- 
    -- CP-element group 363:  transition  input  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	99 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (2) 
      -- CP-element group 363: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_382/SplitProtocol/Update/$exit
      -- CP-element group 363: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_382/SplitProtocol/Update/ca
      -- 
    ca_3769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_382_inst_ack_1, ack => testConfigure_CP_0_elements(363)); -- 
    -- CP-element group 364:  join  transition  output  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	362 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	365 
    -- CP-element group 364:  members (5) 
      -- CP-element group 364: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_379/$exit
      -- CP-element group 364: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/$exit
      -- CP-element group 364: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_382/$exit
      -- CP-element group 364: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_382/SplitProtocol/$exit
      -- CP-element group 364: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_req
      -- 
    phi_stmt_379_req_3770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_379_req_3770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(364), ack => phi_stmt_379_req_0); -- 
    testConfigure_cp_element_group_364: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_364"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(362) & testConfigure_CP_0_elements(363);
      gj_testConfigure_cp_element_group_364 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(364), clk => clk, reset => reset); --
    end block;
    -- CP-element group 365:  join  transition  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	361 
    -- CP-element group 365: 	364 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	373 
    -- CP-element group 365:  members (1) 
      -- CP-element group 365: 	 branch_block_stmt_34/bbx_xnph307_forx_xbody69_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_365: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_365"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(361) & testConfigure_CP_0_elements(364);
      gj_testConfigure_cp_element_group_365 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(365), clk => clk, reset => reset); --
    end block;
    -- CP-element group 366:  transition  input  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	118 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	368 
    -- CP-element group 366:  members (2) 
      -- CP-element group 366: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_372/phi_stmt_372_sources/type_cast_378/SplitProtocol/Sample/$exit
      -- CP-element group 366: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_372/phi_stmt_372_sources/type_cast_378/SplitProtocol/Sample/ra
      -- 
    ra_3790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_378_inst_ack_0, ack => testConfigure_CP_0_elements(366)); -- 
    -- CP-element group 367:  transition  input  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	118 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367:  members (2) 
      -- CP-element group 367: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_372/phi_stmt_372_sources/type_cast_378/SplitProtocol/Update/$exit
      -- CP-element group 367: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_372/phi_stmt_372_sources/type_cast_378/SplitProtocol/Update/ca
      -- 
    ca_3795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_378_inst_ack_1, ack => testConfigure_CP_0_elements(367)); -- 
    -- CP-element group 368:  join  transition  output  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	366 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	372 
    -- CP-element group 368:  members (5) 
      -- CP-element group 368: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_372/$exit
      -- CP-element group 368: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_372/phi_stmt_372_sources/$exit
      -- CP-element group 368: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_372/phi_stmt_372_sources/type_cast_378/$exit
      -- CP-element group 368: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_372/phi_stmt_372_sources/type_cast_378/SplitProtocol/$exit
      -- CP-element group 368: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_372/phi_stmt_372_req
      -- 
    phi_stmt_372_req_3796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_372_req_3796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(368), ack => phi_stmt_372_req_1); -- 
    testConfigure_cp_element_group_368: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_368"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(366) & testConfigure_CP_0_elements(367);
      gj_testConfigure_cp_element_group_368 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(368), clk => clk, reset => reset); --
    end block;
    -- CP-element group 369:  transition  input  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	118 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	371 
    -- CP-element group 369:  members (2) 
      -- CP-element group 369: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_384/SplitProtocol/Sample/$exit
      -- CP-element group 369: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_384/SplitProtocol/Sample/ra
      -- 
    ra_3813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_384_inst_ack_0, ack => testConfigure_CP_0_elements(369)); -- 
    -- CP-element group 370:  transition  input  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	118 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	371 
    -- CP-element group 370:  members (2) 
      -- CP-element group 370: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_384/SplitProtocol/Update/$exit
      -- CP-element group 370: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_384/SplitProtocol/Update/ca
      -- 
    ca_3818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_384_inst_ack_1, ack => testConfigure_CP_0_elements(370)); -- 
    -- CP-element group 371:  join  transition  output  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	369 
    -- CP-element group 371: 	370 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (5) 
      -- CP-element group 371: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_379/$exit
      -- CP-element group 371: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/$exit
      -- CP-element group 371: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_384/$exit
      -- CP-element group 371: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_sources/type_cast_384/SplitProtocol/$exit
      -- CP-element group 371: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/phi_stmt_379/phi_stmt_379_req
      -- 
    phi_stmt_379_req_3819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_379_req_3819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(371), ack => phi_stmt_379_req_1); -- 
    testConfigure_cp_element_group_371: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_371"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(369) & testConfigure_CP_0_elements(370);
      gj_testConfigure_cp_element_group_371 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(371), clk => clk, reset => reset); --
    end block;
    -- CP-element group 372:  join  transition  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	368 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (1) 
      -- CP-element group 372: 	 branch_block_stmt_34/forx_xbody69_forx_xbody69_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_372: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_372"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(368) & testConfigure_CP_0_elements(371);
      gj_testConfigure_cp_element_group_372 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(372), clk => clk, reset => reset); --
    end block;
    -- CP-element group 373:  merge  fork  transition  place  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	365 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373: 	375 
    -- CP-element group 373:  members (2) 
      -- CP-element group 373: 	 branch_block_stmt_34/merge_stmt_371_PhiReqMerge
      -- CP-element group 373: 	 branch_block_stmt_34/merge_stmt_371_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(373) <= OrReduce(testConfigure_CP_0_elements(365) & testConfigure_CP_0_elements(372));
    -- CP-element group 374:  transition  input  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	376 
    -- CP-element group 374:  members (1) 
      -- CP-element group 374: 	 branch_block_stmt_34/merge_stmt_371_PhiAck/phi_stmt_372_ack
      -- 
    phi_stmt_372_ack_3824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_372_ack_0, ack => testConfigure_CP_0_elements(374)); -- 
    -- CP-element group 375:  transition  input  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	373 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	376 
    -- CP-element group 375:  members (1) 
      -- CP-element group 375: 	 branch_block_stmt_34/merge_stmt_371_PhiAck/phi_stmt_379_ack
      -- 
    phi_stmt_379_ack_3825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_379_ack_0, ack => testConfigure_CP_0_elements(375)); -- 
    -- CP-element group 376:  join  fork  transition  place  output  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	374 
    -- CP-element group 376: 	375 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	100 
    -- CP-element group 376: 	101 
    -- CP-element group 376: 	103 
    -- CP-element group 376: 	104 
    -- CP-element group 376: 	107 
    -- CP-element group 376: 	110 
    -- CP-element group 376: 	114 
    -- CP-element group 376:  members (50) 
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/array_obj_ref_388_index_resize_0/$entry
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_update_start_
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/array_obj_ref_388_index_resize_0/$exit
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_402_sample_start_
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/array_obj_ref_388_index_computed_0
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/array_obj_ref_388_index_scaled_0
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/array_obj_ref_388_index_resized_0
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_Update/word_access_complete/word_0/cr
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/array_obj_ref_388_offset_calculated
      -- CP-element group 376: 	 branch_block_stmt_34/merge_stmt_371__exit__
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435__entry__
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/array_obj_ref_388_root_address_calculated
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_Update/word_access_complete/word_0/$entry
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/addr_of_389_update_start_
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/addr_of_389_sample_start_
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_Update/word_access_complete/$entry
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/$entry
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_392_Update/$entry
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_update_start_
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/addr_of_389_complete/req
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/addr_of_389_complete/$entry
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/array_obj_ref_388_final_index_sum_regn/$entry
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/array_obj_ref_388_index_scale_0/scale_rename_ack
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_402_Sample/rr
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/addr_of_389_request/req
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_406_Update/cr
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/addr_of_389_request/$entry
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_422_Update/cr
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_406_Update/$entry
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_422_Update/$entry
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_Update/word_access_complete/word_0/cr
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/array_obj_ref_388_base_plus_offset/sum_rename_ack
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_Update/word_access_complete/word_0/$entry
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_Update/word_access_complete/$entry
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/array_obj_ref_388_base_plus_offset/sum_rename_req
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/ptr_deref_414_Update/$entry
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_406_update_start_
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/type_cast_422_update_start_
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/array_obj_ref_388_base_plus_offset/$exit
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/array_obj_ref_388_base_plus_offset/$entry
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/array_obj_ref_388_final_index_sum_regn/ack
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/array_obj_ref_388_final_index_sum_regn/req
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/array_obj_ref_388_final_index_sum_regn/$exit
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/array_obj_ref_388_index_scale_0/scale_rename_req
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/array_obj_ref_388_index_scale_0/$exit
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/array_obj_ref_388_index_scale_0/$entry
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/array_obj_ref_388_index_resize_0/index_resize_ack
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/array_obj_ref_388_index_resize_0/index_resize_req
      -- CP-element group 376: 	 branch_block_stmt_34/assign_stmt_390_to_assign_stmt_435/RPIPE_ConvTranspose_input_pipe_402_Sample/$entry
      -- CP-element group 376: 	 branch_block_stmt_34/merge_stmt_371_PhiAck/$exit
      -- 
    cr_1195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(376), ack => ptr_deref_392_store_0_req_1); -- 
    req_1145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(376), ack => addr_of_389_final_reg_req_1); -- 
    rr_1204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(376), ack => RPIPE_ConvTranspose_input_pipe_402_inst_req_0); -- 
    req_1140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(376), ack => addr_of_389_final_reg_req_0); -- 
    cr_1223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(376), ack => type_cast_406_inst_req_1); -- 
    cr_1301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(376), ack => type_cast_422_inst_req_1); -- 
    cr_1273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(376), ack => ptr_deref_414_store_0_req_1); -- 
    testConfigure_cp_element_group_376: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_376"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(374) & testConfigure_CP_0_elements(375);
      gj_testConfigure_cp_element_group_376 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(376), clk => clk, reset => reset); --
    end block;
    -- CP-element group 377:  transition  input  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	117 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	379 
    -- CP-element group 377:  members (2) 
      -- CP-element group 377: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_443/phi_stmt_443_sources/type_cast_446/SplitProtocol/Sample/$exit
      -- CP-element group 377: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_443/phi_stmt_443_sources/type_cast_446/SplitProtocol/Sample/ra
      -- 
    ra_3849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_446_inst_ack_0, ack => testConfigure_CP_0_elements(377)); -- 
    -- CP-element group 378:  transition  input  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	117 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	379 
    -- CP-element group 378:  members (2) 
      -- CP-element group 378: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_443/phi_stmt_443_sources/type_cast_446/SplitProtocol/Update/$exit
      -- CP-element group 378: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_443/phi_stmt_443_sources/type_cast_446/SplitProtocol/Update/ca
      -- 
    ca_3854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_446_inst_ack_1, ack => testConfigure_CP_0_elements(378)); -- 
    -- CP-element group 379:  join  transition  output  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	377 
    -- CP-element group 379: 	378 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	383 
    -- CP-element group 379:  members (5) 
      -- CP-element group 379: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_443/$exit
      -- CP-element group 379: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_443/phi_stmt_443_sources/$exit
      -- CP-element group 379: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_443/phi_stmt_443_sources/type_cast_446/$exit
      -- CP-element group 379: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_443/phi_stmt_443_sources/type_cast_446/SplitProtocol/$exit
      -- CP-element group 379: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_443/phi_stmt_443_req
      -- 
    phi_stmt_443_req_3855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_443_req_3855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(379), ack => phi_stmt_443_req_0); -- 
    testConfigure_cp_element_group_379: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_379"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(377) & testConfigure_CP_0_elements(378);
      gj_testConfigure_cp_element_group_379 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(379), clk => clk, reset => reset); --
    end block;
    -- CP-element group 380:  transition  input  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	117 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	382 
    -- CP-element group 380:  members (2) 
      -- CP-element group 380: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_447/phi_stmt_447_sources/type_cast_450/SplitProtocol/Sample/$exit
      -- CP-element group 380: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_447/phi_stmt_447_sources/type_cast_450/SplitProtocol/Sample/ra
      -- 
    ra_3872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_450_inst_ack_0, ack => testConfigure_CP_0_elements(380)); -- 
    -- CP-element group 381:  transition  input  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	117 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	382 
    -- CP-element group 381:  members (2) 
      -- CP-element group 381: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_447/phi_stmt_447_sources/type_cast_450/SplitProtocol/Update/$exit
      -- CP-element group 381: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_447/phi_stmt_447_sources/type_cast_450/SplitProtocol/Update/ca
      -- 
    ca_3877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_450_inst_ack_1, ack => testConfigure_CP_0_elements(381)); -- 
    -- CP-element group 382:  join  transition  output  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	380 
    -- CP-element group 382: 	381 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	383 
    -- CP-element group 382:  members (5) 
      -- CP-element group 382: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_447/$exit
      -- CP-element group 382: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_447/phi_stmt_447_sources/$exit
      -- CP-element group 382: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_447/phi_stmt_447_sources/type_cast_450/$exit
      -- CP-element group 382: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_447/phi_stmt_447_sources/type_cast_450/SplitProtocol/$exit
      -- CP-element group 382: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/phi_stmt_447/phi_stmt_447_req
      -- 
    phi_stmt_447_req_3878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_447_req_3878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(382), ack => phi_stmt_447_req_0); -- 
    testConfigure_cp_element_group_382: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_382"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(380) & testConfigure_CP_0_elements(381);
      gj_testConfigure_cp_element_group_382 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(382), clk => clk, reset => reset); --
    end block;
    -- CP-element group 383:  join  fork  transition  place  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	379 
    -- CP-element group 383: 	382 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	384 
    -- CP-element group 383: 	385 
    -- CP-element group 383:  members (3) 
      -- CP-element group 383: 	 branch_block_stmt_34/forx_xbody69_forx_xend91_PhiReq/$exit
      -- CP-element group 383: 	 branch_block_stmt_34/merge_stmt_442_PhiReqMerge
      -- CP-element group 383: 	 branch_block_stmt_34/merge_stmt_442_PhiAck/$entry
      -- 
    testConfigure_cp_element_group_383: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_383"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(379) & testConfigure_CP_0_elements(382);
      gj_testConfigure_cp_element_group_383 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(383), clk => clk, reset => reset); --
    end block;
    -- CP-element group 384:  transition  input  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	383 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	386 
    -- CP-element group 384:  members (1) 
      -- CP-element group 384: 	 branch_block_stmt_34/merge_stmt_442_PhiAck/phi_stmt_443_ack
      -- 
    phi_stmt_443_ack_3883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_443_ack_0, ack => testConfigure_CP_0_elements(384)); -- 
    -- CP-element group 385:  transition  input  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	383 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	386 
    -- CP-element group 385:  members (1) 
      -- CP-element group 385: 	 branch_block_stmt_34/merge_stmt_442_PhiAck/phi_stmt_447_ack
      -- 
    phi_stmt_447_ack_3884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_447_ack_0, ack => testConfigure_CP_0_elements(385)); -- 
    -- CP-element group 386:  join  transition  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	384 
    -- CP-element group 386: 	385 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	1 
    -- CP-element group 386:  members (1) 
      -- CP-element group 386: 	 branch_block_stmt_34/merge_stmt_442_PhiAck/$exit
      -- 
    testConfigure_cp_element_group_386: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_386"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(384) & testConfigure_CP_0_elements(385);
      gj_testConfigure_cp_element_group_386 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(386), clk => clk, reset => reset); --
    end block;
    -- CP-element group 387:  merge  branch  transition  place  output  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	209 
    -- CP-element group 387: 	254 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	210 
    -- CP-element group 387: 	211 
    -- CP-element group 387:  members (17) 
      -- CP-element group 387: 	 branch_block_stmt_34/merge_stmt_778__exit__
      -- CP-element group 387: 	 branch_block_stmt_34/assign_stmt_784__entry__
      -- CP-element group 387: 	 branch_block_stmt_34/assign_stmt_784__exit__
      -- CP-element group 387: 	 branch_block_stmt_34/if_stmt_785__entry__
      -- CP-element group 387: 	 branch_block_stmt_34/R_cmp211295_786_place
      -- CP-element group 387: 	 branch_block_stmt_34/if_stmt_785_eval_test/$exit
      -- CP-element group 387: 	 branch_block_stmt_34/assign_stmt_784/$exit
      -- CP-element group 387: 	 branch_block_stmt_34/if_stmt_785_eval_test/branch_req
      -- CP-element group 387: 	 branch_block_stmt_34/if_stmt_785_dead_link/$entry
      -- CP-element group 387: 	 branch_block_stmt_34/if_stmt_785_if_link/$entry
      -- CP-element group 387: 	 branch_block_stmt_34/if_stmt_785_else_link/$entry
      -- CP-element group 387: 	 branch_block_stmt_34/assign_stmt_784/$entry
      -- CP-element group 387: 	 branch_block_stmt_34/if_stmt_785_eval_test/$entry
      -- CP-element group 387: 	 branch_block_stmt_34/merge_stmt_778_PhiReqMerge
      -- CP-element group 387: 	 branch_block_stmt_34/merge_stmt_778_PhiAck/$entry
      -- CP-element group 387: 	 branch_block_stmt_34/merge_stmt_778_PhiAck/$exit
      -- CP-element group 387: 	 branch_block_stmt_34/merge_stmt_778_PhiAck/dummy
      -- 
    branch_req_2385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(387), ack => if_stmt_785_branch_req_0); -- 
    testConfigure_CP_0_elements(387) <= OrReduce(testConfigure_CP_0_elements(209) & testConfigure_CP_0_elements(254));
    -- CP-element group 388:  transition  output  delay-element  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	213 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	392 
    -- CP-element group 388:  members (5) 
      -- CP-element group 388: 	 branch_block_stmt_34/bbx_xnph301_forx_xbody153_PhiReq/$exit
      -- CP-element group 388: 	 branch_block_stmt_34/bbx_xnph301_forx_xbody153_PhiReq/phi_stmt_829/$exit
      -- CP-element group 388: 	 branch_block_stmt_34/bbx_xnph301_forx_xbody153_PhiReq/phi_stmt_829/phi_stmt_829_sources/$exit
      -- CP-element group 388: 	 branch_block_stmt_34/bbx_xnph301_forx_xbody153_PhiReq/phi_stmt_829/phi_stmt_829_sources/type_cast_833_konst_delay_trans
      -- CP-element group 388: 	 branch_block_stmt_34/bbx_xnph301_forx_xbody153_PhiReq/phi_stmt_829/phi_stmt_829_req
      -- 
    phi_stmt_829_req_3930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_829_req_3930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(388), ack => phi_stmt_829_req_0); -- 
    -- Element group testConfigure_CP_0_elements(388) is a control-delay.
    cp_element_388_delay: control_delay_element  generic map(name => " 388_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(213), ack => testConfigure_CP_0_elements(388), clk => clk, reset =>reset);
    -- CP-element group 389:  transition  input  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	255 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	391 
    -- CP-element group 389:  members (2) 
      -- CP-element group 389: 	 branch_block_stmt_34/forx_xbody153_forx_xbody153_PhiReq/phi_stmt_829/phi_stmt_829_sources/type_cast_835/SplitProtocol/Sample/$exit
      -- CP-element group 389: 	 branch_block_stmt_34/forx_xbody153_forx_xbody153_PhiReq/phi_stmt_829/phi_stmt_829_sources/type_cast_835/SplitProtocol/Sample/ra
      -- 
    ra_3950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_835_inst_ack_0, ack => testConfigure_CP_0_elements(389)); -- 
    -- CP-element group 390:  transition  input  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	255 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	391 
    -- CP-element group 390:  members (2) 
      -- CP-element group 390: 	 branch_block_stmt_34/forx_xbody153_forx_xbody153_PhiReq/phi_stmt_829/phi_stmt_829_sources/type_cast_835/SplitProtocol/Update/$exit
      -- CP-element group 390: 	 branch_block_stmt_34/forx_xbody153_forx_xbody153_PhiReq/phi_stmt_829/phi_stmt_829_sources/type_cast_835/SplitProtocol/Update/ca
      -- 
    ca_3955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_835_inst_ack_1, ack => testConfigure_CP_0_elements(390)); -- 
    -- CP-element group 391:  join  transition  output  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	389 
    -- CP-element group 391: 	390 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	392 
    -- CP-element group 391:  members (6) 
      -- CP-element group 391: 	 branch_block_stmt_34/forx_xbody153_forx_xbody153_PhiReq/$exit
      -- CP-element group 391: 	 branch_block_stmt_34/forx_xbody153_forx_xbody153_PhiReq/phi_stmt_829/$exit
      -- CP-element group 391: 	 branch_block_stmt_34/forx_xbody153_forx_xbody153_PhiReq/phi_stmt_829/phi_stmt_829_sources/$exit
      -- CP-element group 391: 	 branch_block_stmt_34/forx_xbody153_forx_xbody153_PhiReq/phi_stmt_829/phi_stmt_829_sources/type_cast_835/$exit
      -- CP-element group 391: 	 branch_block_stmt_34/forx_xbody153_forx_xbody153_PhiReq/phi_stmt_829/phi_stmt_829_sources/type_cast_835/SplitProtocol/$exit
      -- CP-element group 391: 	 branch_block_stmt_34/forx_xbody153_forx_xbody153_PhiReq/phi_stmt_829/phi_stmt_829_req
      -- 
    phi_stmt_829_req_3956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_829_req_3956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(391), ack => phi_stmt_829_req_1); -- 
    testConfigure_cp_element_group_391: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_391"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(389) & testConfigure_CP_0_elements(390);
      gj_testConfigure_cp_element_group_391 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(391), clk => clk, reset => reset); --
    end block;
    -- CP-element group 392:  merge  transition  place  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	388 
    -- CP-element group 392: 	391 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	393 
    -- CP-element group 392:  members (2) 
      -- CP-element group 392: 	 branch_block_stmt_34/merge_stmt_828_PhiReqMerge
      -- CP-element group 392: 	 branch_block_stmt_34/merge_stmt_828_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(392) <= OrReduce(testConfigure_CP_0_elements(388) & testConfigure_CP_0_elements(391));
    -- CP-element group 393:  fork  transition  place  input  output  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	392 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	214 
    -- CP-element group 393: 	215 
    -- CP-element group 393: 	217 
    -- CP-element group 393: 	218 
    -- CP-element group 393: 	221 
    -- CP-element group 393: 	225 
    -- CP-element group 393: 	229 
    -- CP-element group 393: 	233 
    -- CP-element group 393: 	237 
    -- CP-element group 393: 	241 
    -- CP-element group 393: 	245 
    -- CP-element group 393: 	249 
    -- CP-element group 393: 	252 
    -- CP-element group 393:  members (56) 
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_final_index_sum_regn_Sample/req
      -- CP-element group 393: 	 branch_block_stmt_34/merge_stmt_828__exit__
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991__entry__
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_final_index_sum_regn_Update/req
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_final_index_sum_regn_Update/$entry
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_index_resize_1/$exit
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_862_update_start_
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_898_update_start_
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_862_Update/$entry
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_849_update_start_
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/$entry
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_862_Update/cr
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/addr_of_842_update_start_
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_index_resized_1
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_index_scaled_1
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_index_computed_1
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_index_resize_1/$entry
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_916_Update/cr
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_845_Sample/rr
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_final_index_sum_regn_Sample/$entry
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_845_Sample/$entry
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_898_Update/cr
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_880_update_start_
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_916_Update/$entry
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_final_index_sum_regn_update_start
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/RPIPE_ConvTranspose_input_pipe_845_sample_start_
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_index_scale_1/scale_rename_ack
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_index_scale_1/scale_rename_req
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_index_scale_1/$exit
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_880_Update/cr
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/addr_of_842_complete/req
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_index_scale_1/$entry
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_index_resize_1/index_resize_ack
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/addr_of_842_complete/$entry
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_916_update_start_
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_849_Update/cr
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_849_Update/$entry
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_880_Update/$entry
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/array_obj_ref_841_index_resize_1/index_resize_req
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_898_Update/$entry
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_934_update_start_
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_934_Update/$entry
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_934_Update/cr
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_952_update_start_
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_952_Update/$entry
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_952_Update/cr
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_970_update_start_
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_970_Update/$entry
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/type_cast_970_Update/cr
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_update_start_
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_Update/$entry
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_Update/word_access_complete/$entry
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_Update/word_access_complete/word_0/$entry
      -- CP-element group 393: 	 branch_block_stmt_34/assign_stmt_843_to_assign_stmt_991/ptr_deref_978_Update/word_access_complete/word_0/cr
      -- CP-element group 393: 	 branch_block_stmt_34/merge_stmt_828_PhiAck/$exit
      -- CP-element group 393: 	 branch_block_stmt_34/merge_stmt_828_PhiAck/phi_stmt_829_ack
      -- 
    phi_stmt_829_ack_3961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_829_ack_0, ack => testConfigure_CP_0_elements(393)); -- 
    req_2441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(393), ack => array_obj_ref_841_index_offset_req_0); -- 
    req_2446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(393), ack => array_obj_ref_841_index_offset_req_1); -- 
    cr_2517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(393), ack => type_cast_862_inst_req_1); -- 
    cr_2601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(393), ack => type_cast_916_inst_req_1); -- 
    rr_2470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(393), ack => RPIPE_ConvTranspose_input_pipe_845_inst_req_0); -- 
    cr_2573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(393), ack => type_cast_898_inst_req_1); -- 
    cr_2545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(393), ack => type_cast_880_inst_req_1); -- 
    req_2461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(393), ack => addr_of_842_final_reg_req_1); -- 
    cr_2489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(393), ack => type_cast_849_inst_req_1); -- 
    cr_2629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(393), ack => type_cast_934_inst_req_1); -- 
    cr_2657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(393), ack => type_cast_952_inst_req_1); -- 
    cr_2685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(393), ack => type_cast_970_inst_req_1); -- 
    cr_2735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(393), ack => ptr_deref_978_store_0_req_1); -- 
    -- CP-element group 394:  transition  output  delay-element  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	257 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	398 
    -- CP-element group 394:  members (5) 
      -- CP-element group 394: 	 branch_block_stmt_34/bbx_xnph297_forx_xbody213_PhiReq/$exit
      -- CP-element group 394: 	 branch_block_stmt_34/bbx_xnph297_forx_xbody213_PhiReq/phi_stmt_1036/$exit
      -- CP-element group 394: 	 branch_block_stmt_34/bbx_xnph297_forx_xbody213_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/$exit
      -- CP-element group 394: 	 branch_block_stmt_34/bbx_xnph297_forx_xbody213_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1040_konst_delay_trans
      -- CP-element group 394: 	 branch_block_stmt_34/bbx_xnph297_forx_xbody213_PhiReq/phi_stmt_1036/phi_stmt_1036_req
      -- 
    phi_stmt_1036_req_3984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1036_req_3984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(394), ack => phi_stmt_1036_req_0); -- 
    -- Element group testConfigure_CP_0_elements(394) is a control-delay.
    cp_element_394_delay: control_delay_element  generic map(name => " 394_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(257), ack => testConfigure_CP_0_elements(394), clk => clk, reset =>reset);
    -- CP-element group 395:  transition  input  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	299 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	397 
    -- CP-element group 395:  members (2) 
      -- CP-element group 395: 	 branch_block_stmt_34/forx_xbody213_forx_xbody213_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/SplitProtocol/Sample/$exit
      -- CP-element group 395: 	 branch_block_stmt_34/forx_xbody213_forx_xbody213_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/SplitProtocol/Sample/ra
      -- 
    ra_4004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1042_inst_ack_0, ack => testConfigure_CP_0_elements(395)); -- 
    -- CP-element group 396:  transition  input  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	299 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	397 
    -- CP-element group 396:  members (2) 
      -- CP-element group 396: 	 branch_block_stmt_34/forx_xbody213_forx_xbody213_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/SplitProtocol/Update/$exit
      -- CP-element group 396: 	 branch_block_stmt_34/forx_xbody213_forx_xbody213_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/SplitProtocol/Update/ca
      -- 
    ca_4009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1042_inst_ack_1, ack => testConfigure_CP_0_elements(396)); -- 
    -- CP-element group 397:  join  transition  output  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	395 
    -- CP-element group 397: 	396 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	398 
    -- CP-element group 397:  members (6) 
      -- CP-element group 397: 	 branch_block_stmt_34/forx_xbody213_forx_xbody213_PhiReq/$exit
      -- CP-element group 397: 	 branch_block_stmt_34/forx_xbody213_forx_xbody213_PhiReq/phi_stmt_1036/$exit
      -- CP-element group 397: 	 branch_block_stmt_34/forx_xbody213_forx_xbody213_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/$exit
      -- CP-element group 397: 	 branch_block_stmt_34/forx_xbody213_forx_xbody213_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/$exit
      -- CP-element group 397: 	 branch_block_stmt_34/forx_xbody213_forx_xbody213_PhiReq/phi_stmt_1036/phi_stmt_1036_sources/type_cast_1042/SplitProtocol/$exit
      -- CP-element group 397: 	 branch_block_stmt_34/forx_xbody213_forx_xbody213_PhiReq/phi_stmt_1036/phi_stmt_1036_req
      -- 
    phi_stmt_1036_req_4010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1036_req_4010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(397), ack => phi_stmt_1036_req_1); -- 
    testConfigure_cp_element_group_397: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_397"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(395) & testConfigure_CP_0_elements(396);
      gj_testConfigure_cp_element_group_397 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(397), clk => clk, reset => reset); --
    end block;
    -- CP-element group 398:  merge  transition  place  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	394 
    -- CP-element group 398: 	397 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	399 
    -- CP-element group 398:  members (2) 
      -- CP-element group 398: 	 branch_block_stmt_34/merge_stmt_1035_PhiReqMerge
      -- CP-element group 398: 	 branch_block_stmt_34/merge_stmt_1035_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(398) <= OrReduce(testConfigure_CP_0_elements(394) & testConfigure_CP_0_elements(397));
    -- CP-element group 399:  fork  transition  place  input  output  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	398 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	258 
    -- CP-element group 399: 	259 
    -- CP-element group 399: 	261 
    -- CP-element group 399: 	262 
    -- CP-element group 399: 	265 
    -- CP-element group 399: 	269 
    -- CP-element group 399: 	273 
    -- CP-element group 399: 	277 
    -- CP-element group 399: 	281 
    -- CP-element group 399: 	285 
    -- CP-element group 399: 	289 
    -- CP-element group 399: 	293 
    -- CP-element group 399: 	296 
    -- CP-element group 399:  members (56) 
      -- CP-element group 399: 	 branch_block_stmt_34/merge_stmt_1035__exit__
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198__entry__
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/$entry
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/addr_of_1049_update_start_
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_index_resized_1
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_index_scaled_1
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_index_computed_1
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_index_resize_1/$entry
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_index_resize_1/$exit
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_index_resize_1/index_resize_req
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_index_resize_1/index_resize_ack
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_index_scale_1/$entry
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_index_scale_1/$exit
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_index_scale_1/scale_rename_req
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_index_scale_1/scale_rename_ack
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_final_index_sum_regn_update_start
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_final_index_sum_regn_Sample/$entry
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_final_index_sum_regn_Sample/req
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_final_index_sum_regn_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/array_obj_ref_1048_final_index_sum_regn_Update/req
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/addr_of_1049_complete/$entry
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/addr_of_1049_complete/req
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1052_sample_start_
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1052_Sample/$entry
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/RPIPE_ConvTranspose_input_pipe_1052_Sample/rr
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1056_update_start_
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1056_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1056_Update/cr
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1069_update_start_
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1069_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1069_Update/cr
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1087_update_start_
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1087_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1087_Update/cr
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1105_update_start_
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1105_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1105_Update/cr
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1123_update_start_
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1123_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1123_Update/cr
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1141_update_start_
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1141_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1141_Update/cr
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1159_update_start_
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1159_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1159_Update/cr
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1177_update_start_
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1177_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/type_cast_1177_Update/cr
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_update_start_
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_Update/word_access_complete/$entry
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_Update/word_access_complete/word_0/$entry
      -- CP-element group 399: 	 branch_block_stmt_34/assign_stmt_1050_to_assign_stmt_1198/ptr_deref_1185_Update/word_access_complete/word_0/cr
      -- CP-element group 399: 	 branch_block_stmt_34/merge_stmt_1035_PhiAck/$exit
      -- CP-element group 399: 	 branch_block_stmt_34/merge_stmt_1035_PhiAck/phi_stmt_1036_ack
      -- 
    phi_stmt_1036_ack_4015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1036_ack_0, ack => testConfigure_CP_0_elements(399)); -- 
    req_2800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(399), ack => array_obj_ref_1048_index_offset_req_0); -- 
    req_2805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(399), ack => array_obj_ref_1048_index_offset_req_1); -- 
    req_2820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(399), ack => addr_of_1049_final_reg_req_1); -- 
    rr_2829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(399), ack => RPIPE_ConvTranspose_input_pipe_1052_inst_req_0); -- 
    cr_2848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(399), ack => type_cast_1056_inst_req_1); -- 
    cr_2876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(399), ack => type_cast_1069_inst_req_1); -- 
    cr_2904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(399), ack => type_cast_1087_inst_req_1); -- 
    cr_2932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(399), ack => type_cast_1105_inst_req_1); -- 
    cr_2960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(399), ack => type_cast_1123_inst_req_1); -- 
    cr_2988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(399), ack => type_cast_1141_inst_req_1); -- 
    cr_3016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(399), ack => type_cast_1159_inst_req_1); -- 
    cr_3044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(399), ack => type_cast_1177_inst_req_1); -- 
    cr_3094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(399), ack => ptr_deref_1185_store_0_req_1); -- 
    -- CP-element group 400:  merge  place  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	211 
    -- CP-element group 400: 	298 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	401 
    -- CP-element group 400:  members (1) 
      -- CP-element group 400: 	 branch_block_stmt_34/merge_stmt_1207_PhiReqMerge
      -- 
    testConfigure_CP_0_elements(400) <= OrReduce(testConfigure_CP_0_elements(211) & testConfigure_CP_0_elements(298));
    -- CP-element group 401:  join  fork  transition  place  output  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	400 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	300 
    -- CP-element group 401: 	301 
    -- CP-element group 401: 	303 
    -- CP-element group 401: 	304 
    -- CP-element group 401: 	305 
    -- CP-element group 401: 	307 
    -- CP-element group 401: 	308 
    -- CP-element group 401: 	309 
    -- CP-element group 401: 	311 
    -- CP-element group 401:  members (93) 
      -- CP-element group 401: 	 branch_block_stmt_34/merge_stmt_1207__exit__
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271__entry__
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_base_addr_resize/base_resize_req
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_Update/word_access_complete/word_0/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_base_plus_offset/sum_rename_req
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_word_address_calculated
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_base_address_calculated
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_root_address_calculated
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_base_addr_resize/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_root_address_calculated
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_base_address_resized
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_base_address_calculated
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_base_plus_offset/sum_rename_ack
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1222_update_start_
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_update_start_
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_base_addr_resize/base_resize_ack
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_base_addr_resize/$exit
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1222_Update/cr
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_base_address_resized
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_base_plus_offset/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_base_plus_offset/$exit
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_base_addr_resize/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_word_address_calculated
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1222_Update/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_root_address_calculated
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_base_addr_resize/base_resize_ack
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_word_address_calculated
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_sample_start_
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_word_addrgen/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_word_addrgen/$exit
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_base_address_resized
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_base_addr_resize/$exit
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_Update/word_access_complete/word_0/cr
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_word_addrgen/root_register_req
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_word_addrgen/root_register_ack
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_base_addr_resize/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_base_addr_resize/$exit
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_base_addr_resize/base_resize_req
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_Sample/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_sample_start_
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1238_Update/cr
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_Update/word_access_complete/word_0/cr
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1238_Update/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_base_address_calculated
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_Update/word_access_complete/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_update_start_
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1238_update_start_
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_update_start_
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_Update/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_sample_start_
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_Sample/word_access_start/word_0/rr
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_Sample/word_access_start/word_0/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1250_Sample/word_access_start/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_Update/word_access_complete/word_0/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_Update/word_access_complete/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_Update/word_access_complete/word_0/cr
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_Update/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_Update/word_access_complete/word_0/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_Sample/word_access_start/word_0/rr
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_Update/word_access_complete/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_Sample/word_access_start/word_0/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_Update/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1254_Update/cr
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_Sample/word_access_start/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_Sample/word_access_start/word_0/rr
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1254_Update/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_Sample/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_Sample/word_access_start/word_0/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_Sample/word_access_start/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_Sample/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_word_addrgen/root_register_ack
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_word_addrgen/root_register_req
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/type_cast_1254_update_start_
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_word_addrgen/$exit
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_word_addrgen/root_register_ack
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_word_addrgen/root_register_req
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_word_addrgen/$exit
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_word_addrgen/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_base_plus_offset/sum_rename_ack
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_word_addrgen/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_base_plus_offset/sum_rename_ack
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_base_plus_offset/sum_rename_req
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_base_plus_offset/sum_rename_req
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_base_plus_offset/$exit
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_base_plus_offset/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_base_addr_resize/base_resize_ack
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1234_base_addr_resize/base_resize_req
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_base_plus_offset/$exit
      -- CP-element group 401: 	 branch_block_stmt_34/assign_stmt_1215_to_assign_stmt_1271/ptr_deref_1218_base_plus_offset/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/merge_stmt_1207_PhiAck/$entry
      -- CP-element group 401: 	 branch_block_stmt_34/merge_stmt_1207_PhiAck/$exit
      -- CP-element group 401: 	 branch_block_stmt_34/merge_stmt_1207_PhiAck/dummy
      -- 
    cr_3180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(401), ack => type_cast_1222_inst_req_1); -- 
    cr_3289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(401), ack => ptr_deref_1250_load_0_req_1); -- 
    cr_3244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(401), ack => type_cast_1238_inst_req_1); -- 
    cr_3161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(401), ack => ptr_deref_1218_load_0_req_1); -- 
    rr_3278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(401), ack => ptr_deref_1250_load_0_req_0); -- 
    cr_3225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(401), ack => ptr_deref_1234_load_0_req_1); -- 
    rr_3150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(401), ack => ptr_deref_1218_load_0_req_0); -- 
    cr_3308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(401), ack => type_cast_1254_inst_req_1); -- 
    rr_3214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(401), ack => ptr_deref_1234_load_0_req_0); -- 
    testConfigure_CP_0_elements(401) <= testConfigure_CP_0_elements(400);
    -- CP-element group 402:  transition  output  delay-element  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	316 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	406 
    -- CP-element group 402:  members (5) 
      -- CP-element group 402: 	 branch_block_stmt_34/bbx_xnph_forx_xbody283_PhiReq/$exit
      -- CP-element group 402: 	 branch_block_stmt_34/bbx_xnph_forx_xbody283_PhiReq/phi_stmt_1316/$exit
      -- CP-element group 402: 	 branch_block_stmt_34/bbx_xnph_forx_xbody283_PhiReq/phi_stmt_1316/phi_stmt_1316_sources/$exit
      -- CP-element group 402: 	 branch_block_stmt_34/bbx_xnph_forx_xbody283_PhiReq/phi_stmt_1316/phi_stmt_1316_sources/type_cast_1320_konst_delay_trans
      -- CP-element group 402: 	 branch_block_stmt_34/bbx_xnph_forx_xbody283_PhiReq/phi_stmt_1316/phi_stmt_1316_req
      -- 
    phi_stmt_1316_req_4061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1316_req_4061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(402), ack => phi_stmt_1316_req_0); -- 
    -- Element group testConfigure_CP_0_elements(402) is a control-delay.
    cp_element_402_delay: control_delay_element  generic map(name => " 402_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(316), ack => testConfigure_CP_0_elements(402), clk => clk, reset =>reset);
    -- CP-element group 403:  transition  input  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	325 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	405 
    -- CP-element group 403:  members (2) 
      -- CP-element group 403: 	 branch_block_stmt_34/forx_xbody283_forx_xbody283_PhiReq/phi_stmt_1316/phi_stmt_1316_sources/type_cast_1322/SplitProtocol/Sample/$exit
      -- CP-element group 403: 	 branch_block_stmt_34/forx_xbody283_forx_xbody283_PhiReq/phi_stmt_1316/phi_stmt_1316_sources/type_cast_1322/SplitProtocol/Sample/ra
      -- 
    ra_4081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1322_inst_ack_0, ack => testConfigure_CP_0_elements(403)); -- 
    -- CP-element group 404:  transition  input  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	325 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	405 
    -- CP-element group 404:  members (2) 
      -- CP-element group 404: 	 branch_block_stmt_34/forx_xbody283_forx_xbody283_PhiReq/phi_stmt_1316/phi_stmt_1316_sources/type_cast_1322/SplitProtocol/Update/$exit
      -- CP-element group 404: 	 branch_block_stmt_34/forx_xbody283_forx_xbody283_PhiReq/phi_stmt_1316/phi_stmt_1316_sources/type_cast_1322/SplitProtocol/Update/ca
      -- 
    ca_4086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1322_inst_ack_1, ack => testConfigure_CP_0_elements(404)); -- 
    -- CP-element group 405:  join  transition  output  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	403 
    -- CP-element group 405: 	404 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	406 
    -- CP-element group 405:  members (6) 
      -- CP-element group 405: 	 branch_block_stmt_34/forx_xbody283_forx_xbody283_PhiReq/$exit
      -- CP-element group 405: 	 branch_block_stmt_34/forx_xbody283_forx_xbody283_PhiReq/phi_stmt_1316/$exit
      -- CP-element group 405: 	 branch_block_stmt_34/forx_xbody283_forx_xbody283_PhiReq/phi_stmt_1316/phi_stmt_1316_sources/$exit
      -- CP-element group 405: 	 branch_block_stmt_34/forx_xbody283_forx_xbody283_PhiReq/phi_stmt_1316/phi_stmt_1316_sources/type_cast_1322/$exit
      -- CP-element group 405: 	 branch_block_stmt_34/forx_xbody283_forx_xbody283_PhiReq/phi_stmt_1316/phi_stmt_1316_sources/type_cast_1322/SplitProtocol/$exit
      -- CP-element group 405: 	 branch_block_stmt_34/forx_xbody283_forx_xbody283_PhiReq/phi_stmt_1316/phi_stmt_1316_req
      -- 
    phi_stmt_1316_req_4087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1316_req_4087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(405), ack => phi_stmt_1316_req_1); -- 
    testConfigure_cp_element_group_405: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_405"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(403) & testConfigure_CP_0_elements(404);
      gj_testConfigure_cp_element_group_405 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(405), clk => clk, reset => reset); --
    end block;
    -- CP-element group 406:  merge  transition  place  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	402 
    -- CP-element group 406: 	405 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	407 
    -- CP-element group 406:  members (2) 
      -- CP-element group 406: 	 branch_block_stmt_34/merge_stmt_1315_PhiReqMerge
      -- CP-element group 406: 	 branch_block_stmt_34/merge_stmt_1315_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(406) <= OrReduce(testConfigure_CP_0_elements(402) & testConfigure_CP_0_elements(405));
    -- CP-element group 407:  fork  transition  place  input  output  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	406 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	317 
    -- CP-element group 407: 	318 
    -- CP-element group 407: 	320 
    -- CP-element group 407: 	322 
    -- CP-element group 407:  members (29) 
      -- CP-element group 407: 	 branch_block_stmt_34/merge_stmt_1315__exit__
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346__entry__
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_index_scale_1/scale_rename_ack
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_index_resize_1/index_resize_ack
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_index_scale_1/$exit
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_Update/word_access_complete/word_0/cr
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_index_scale_1/scale_rename_req
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_index_resize_1/index_resize_req
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_final_index_sum_regn_update_start
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_final_index_sum_regn_Sample/$entry
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_final_index_sum_regn_Sample/req
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_Update/word_access_complete/word_0/$entry
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_index_scale_1/$entry
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_final_index_sum_regn_Update/$entry
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_Update/word_access_complete/$entry
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_final_index_sum_regn_Update/req
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_index_resize_1/$exit
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_index_resize_1/$entry
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_Update/$entry
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_index_computed_1
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_index_scaled_1
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/array_obj_ref_1328_index_resized_1
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/addr_of_1329_update_start_
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/$entry
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/ptr_deref_1332_update_start_
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/addr_of_1329_complete/req
      -- CP-element group 407: 	 branch_block_stmt_34/assign_stmt_1330_to_assign_stmt_1346/addr_of_1329_complete/$entry
      -- CP-element group 407: 	 branch_block_stmt_34/merge_stmt_1315_PhiAck/$exit
      -- CP-element group 407: 	 branch_block_stmt_34/merge_stmt_1315_PhiAck/phi_stmt_1316_ack
      -- 
    phi_stmt_1316_ack_4092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1316_ack_0, ack => testConfigure_CP_0_elements(407)); -- 
    cr_3443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(407), ack => ptr_deref_1332_store_0_req_1); -- 
    req_3373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(407), ack => array_obj_ref_1328_index_offset_req_0); -- 
    req_3378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(407), ack => array_obj_ref_1328_index_offset_req_1); -- 
    req_3393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(407), ack => addr_of_1329_final_reg_req_1); -- 
    -- CP-element group 408:  merge  transition  place  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	314 
    -- CP-element group 408: 	324 
    -- CP-element group 408: successors 
    -- CP-element group 408:  members (20) 
      -- CP-element group 408: 	 $exit
      -- CP-element group 408: 	 branch_block_stmt_34/$exit
      -- CP-element group 408: 	 branch_block_stmt_34/branch_block_stmt_34__exit__
      -- CP-element group 408: 	 branch_block_stmt_34/merge_stmt_1355__exit__
      -- CP-element group 408: 	 branch_block_stmt_34/assign_stmt_1359__entry__
      -- CP-element group 408: 	 branch_block_stmt_34/assign_stmt_1359__exit__
      -- CP-element group 408: 	 branch_block_stmt_34/return__
      -- CP-element group 408: 	 branch_block_stmt_34/merge_stmt_1361__exit__
      -- CP-element group 408: 	 branch_block_stmt_34/assign_stmt_1359/$entry
      -- CP-element group 408: 	 branch_block_stmt_34/assign_stmt_1359/$exit
      -- CP-element group 408: 	 branch_block_stmt_34/merge_stmt_1355_PhiReqMerge
      -- CP-element group 408: 	 branch_block_stmt_34/merge_stmt_1355_PhiAck/$entry
      -- CP-element group 408: 	 branch_block_stmt_34/merge_stmt_1355_PhiAck/$exit
      -- CP-element group 408: 	 branch_block_stmt_34/merge_stmt_1355_PhiAck/dummy
      -- CP-element group 408: 	 branch_block_stmt_34/return___PhiReq/$entry
      -- CP-element group 408: 	 branch_block_stmt_34/return___PhiReq/$exit
      -- CP-element group 408: 	 branch_block_stmt_34/merge_stmt_1361_PhiReqMerge
      -- CP-element group 408: 	 branch_block_stmt_34/merge_stmt_1361_PhiAck/$entry
      -- CP-element group 408: 	 branch_block_stmt_34/merge_stmt_1361_PhiAck/$exit
      -- CP-element group 408: 	 branch_block_stmt_34/merge_stmt_1361_PhiAck/dummy
      -- 
    testConfigure_CP_0_elements(408) <= OrReduce(testConfigure_CP_0_elements(314) & testConfigure_CP_0_elements(324));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar332_1047_resized : std_logic_vector(10 downto 0);
    signal R_indvar332_1047_scaled : std_logic_vector(10 downto 0);
    signal R_indvar348_840_resized : std_logic_vector(13 downto 0);
    signal R_indvar348_840_scaled : std_logic_vector(13 downto 0);
    signal R_indvar364_387_resized : std_logic_vector(0 downto 0);
    signal R_indvar364_387_scaled : std_logic_vector(0 downto 0);
    signal R_indvar367_290_resized : std_logic_vector(6 downto 0);
    signal R_indvar367_290_scaled : std_logic_vector(6 downto 0);
    signal R_indvar372_130_resized : std_logic_vector(6 downto 0);
    signal R_indvar372_130_scaled : std_logic_vector(6 downto 0);
    signal R_indvar_1327_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1327_scaled : std_logic_vector(13 downto 0);
    signal STORE_padding_452_data_0 : std_logic_vector(15 downto 0);
    signal STORE_padding_452_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_padding_477_data_0 : std_logic_vector(15 downto 0);
    signal STORE_padding_477_word_address_0 : std_logic_vector(0 downto 0);
    signal add108_516 : std_logic_vector(15 downto 0);
    signal add117_565 : std_logic_vector(15 downto 0);
    signal add126_614 : std_logic_vector(15 downto 0);
    signal add162_868 : std_logic_vector(63 downto 0);
    signal add168_886 : std_logic_vector(63 downto 0);
    signal add174_904 : std_logic_vector(63 downto 0);
    signal add180_922 : std_logic_vector(63 downto 0);
    signal add186_940 : std_logic_vector(63 downto 0);
    signal add192_958 : std_logic_vector(63 downto 0);
    signal add198_976 : std_logic_vector(63 downto 0);
    signal add21_155 : std_logic_vector(15 downto 0);
    signal add223_1075 : std_logic_vector(63 downto 0);
    signal add229_1093 : std_logic_vector(63 downto 0);
    signal add235_1111 : std_logic_vector(63 downto 0);
    signal add241_1129 : std_logic_vector(63 downto 0);
    signal add247_1147 : std_logic_vector(63 downto 0);
    signal add253_1165 : std_logic_vector(63 downto 0);
    signal add259_1183 : std_logic_vector(63 downto 0);
    signal add34_243 : std_logic_vector(15 downto 0);
    signal add56_322 : std_logic_vector(15 downto 0);
    signal add83_412 : std_logic_vector(15 downto 0);
    signal add99_476 : std_logic_vector(15 downto 0);
    signal add_69 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1048_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1048_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1048_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1048_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1048_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1048_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_131_constant_part_of_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_131_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_131_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_131_offset_scale_factor_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_131_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_131_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_1328_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1328_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1328_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1328_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1328_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1328_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_291_constant_part_of_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_291_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_291_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_291_offset_scale_factor_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_291_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_291_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_388_final_offset : std_logic_vector(0 downto 0);
    signal array_obj_ref_388_offset_scale_factor_0 : std_logic_vector(0 downto 0);
    signal array_obj_ref_388_resized_base_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_388_root_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_841_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_841_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_841_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_841_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_841_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_841_root_address : std_logic_vector(13 downto 0);
    signal arrayidx202_843 : std_logic_vector(31 downto 0);
    signal arrayidx25_133 : std_logic_vector(31 downto 0);
    signal arrayidx263_1050 : std_logic_vector(31 downto 0);
    signal arrayidx286_1330 : std_logic_vector(31 downto 0);
    signal arrayidx60_293 : std_logic_vector(31 downto 0);
    signal arrayidx87_390 : std_logic_vector(31 downto 0);
    signal call101_482 : std_logic_vector(7 downto 0);
    signal call10317_89 : std_logic_vector(7 downto 0);
    signal call106_507 : std_logic_vector(7 downto 0);
    signal call10_190 : std_logic_vector(7 downto 0);
    signal call110_531 : std_logic_vector(7 downto 0);
    signal call115_556 : std_logic_vector(7 downto 0);
    signal call119_580 : std_logic_vector(7 downto 0);
    signal call124_605 : std_logic_vector(7 downto 0);
    signal call155_846 : std_logic_vector(7 downto 0);
    signal call159_859 : std_logic_vector(7 downto 0);
    signal call165_877 : std_logic_vector(7 downto 0);
    signal call171_895 : std_logic_vector(7 downto 0);
    signal call177_913 : std_logic_vector(7 downto 0);
    signal call183_931 : std_logic_vector(7 downto 0);
    signal call189_949 : std_logic_vector(7 downto 0);
    signal call195_967 : std_logic_vector(7 downto 0);
    signal call19_146 : std_logic_vector(7 downto 0);
    signal call216_1053 : std_logic_vector(7 downto 0);
    signal call220_1066 : std_logic_vector(7 downto 0);
    signal call226_1084 : std_logic_vector(7 downto 0);
    signal call232_1102 : std_logic_vector(7 downto 0);
    signal call238_1120 : std_logic_vector(7 downto 0);
    signal call244_1138 : std_logic_vector(7 downto 0);
    signal call250_1156 : std_logic_vector(7 downto 0);
    signal call256_1174 : std_logic_vector(7 downto 0);
    signal call2_60 : std_logic_vector(7 downto 0);
    signal call32_234 : std_logic_vector(7 downto 0);
    signal call43_296 : std_logic_vector(7 downto 0);
    signal call54_313 : std_logic_vector(7 downto 0);
    signal call70303_365 : std_logic_vector(7 downto 0);
    signal call70_419 : std_logic_vector(7 downto 0);
    signal call70x_xlcssa_447 : std_logic_vector(7 downto 0);
    signal call81_403 : std_logic_vector(7 downto 0);
    signal call97_467 : std_logic_vector(7 downto 0);
    signal call_37 : std_logic_vector(7 downto 0);
    signal cmp151299_769 : std_logic_vector(0 downto 0);
    signal cmp211295_784 : std_logic_vector(0 downto 0);
    signal cmp281292_1271 : std_logic_vector(0 downto 0);
    signal cmp316_86 : std_logic_vector(0 downto 0);
    signal cmp40311_259 : std_logic_vector(0 downto 0);
    signal cmp40_353 : std_logic_vector(0 downto 0);
    signal cmp_187 : std_logic_vector(0 downto 0);
    signal conv102_486 : std_logic_vector(15 downto 0);
    signal conv107_511 : std_logic_vector(15 downto 0);
    signal conv111_535 : std_logic_vector(15 downto 0);
    signal conv11318_93 : std_logic_vector(15 downto 0);
    signal conv11320_110 : std_logic_vector(15 downto 0);
    signal conv116_560 : std_logic_vector(15 downto 0);
    signal conv11_194 : std_logic_vector(15 downto 0);
    signal conv11x_xlcssa1_202 : std_logic_vector(15 downto 0);
    signal conv11x_xlcssa_209 : std_logic_vector(15 downto 0);
    signal conv120_584 : std_logic_vector(15 downto 0);
    signal conv125_609 : std_logic_vector(15 downto 0);
    signal conv130_642 : std_logic_vector(31 downto 0);
    signal conv132_658 : std_logic_vector(31 downto 0);
    signal conv134_674 : std_logic_vector(31 downto 0);
    signal conv138_700 : std_logic_vector(31 downto 0);
    signal conv140_716 : std_logic_vector(31 downto 0);
    signal conv143_732 : std_logic_vector(31 downto 0);
    signal conv146_748 : std_logic_vector(31 downto 0);
    signal conv156_850 : std_logic_vector(63 downto 0);
    signal conv161_863 : std_logic_vector(63 downto 0);
    signal conv167_881 : std_logic_vector(63 downto 0);
    signal conv173_899 : std_logic_vector(63 downto 0);
    signal conv179_917 : std_logic_vector(63 downto 0);
    signal conv185_935 : std_logic_vector(63 downto 0);
    signal conv191_953 : std_logic_vector(63 downto 0);
    signal conv197_971 : std_logic_vector(63 downto 0);
    signal conv20_150 : std_logic_vector(15 downto 0);
    signal conv217_1057 : std_logic_vector(63 downto 0);
    signal conv222_1070 : std_logic_vector(63 downto 0);
    signal conv228_1088 : std_logic_vector(63 downto 0);
    signal conv234_1106 : std_logic_vector(63 downto 0);
    signal conv240_1124 : std_logic_vector(63 downto 0);
    signal conv246_1142 : std_logic_vector(63 downto 0);
    signal conv252_1160 : std_logic_vector(63 downto 0);
    signal conv258_1178 : std_logic_vector(63 downto 0);
    signal conv270_1223 : std_logic_vector(31 downto 0);
    signal conv272_1239 : std_logic_vector(31 downto 0);
    signal conv275_1255 : std_logic_vector(31 downto 0);
    signal conv33_238 : std_logic_vector(15 downto 0);
    signal conv39_346 : std_logic_vector(31 downto 0);
    signal conv3_64 : std_logic_vector(15 downto 0);
    signal conv44_300 : std_logic_vector(15 downto 0);
    signal conv55_317 : std_logic_vector(15 downto 0);
    signal conv71304_369 : std_logic_vector(15 downto 0);
    signal conv71306_379 : std_logic_vector(15 downto 0);
    signal conv71_423 : std_logic_vector(15 downto 0);
    signal conv71x_xlcssa_443 : std_logic_vector(15 downto 0);
    signal conv82_407 : std_logic_vector(15 downto 0);
    signal conv8_179 : std_logic_vector(31 downto 0);
    signal conv95_458 : std_logic_vector(15 downto 0);
    signal conv98_471 : std_logic_vector(15 downto 0);
    signal conv_41 : std_logic_vector(15 downto 0);
    signal exitcond5_1346 : std_logic_vector(0 downto 0);
    signal exitcond6_991 : std_logic_vector(0 downto 0);
    signal exitcond7_435 : std_logic_vector(0 downto 0);
    signal exitcond_1198 : std_logic_vector(0 downto 0);
    signal iNsTr_11_249 : std_logic_vector(31 downto 0);
    signal iNsTr_1_47 : std_logic_vector(31 downto 0);
    signal iNsTr_21_171 : std_logic_vector(31 downto 0);
    signal iNsTr_33_338 : std_logic_vector(31 downto 0);
    signal iNsTr_40_494 : std_logic_vector(31 downto 0);
    signal iNsTr_43_524 : std_logic_vector(31 downto 0);
    signal iNsTr_46_543 : std_logic_vector(31 downto 0);
    signal iNsTr_49_573 : std_logic_vector(31 downto 0);
    signal iNsTr_4_75 : std_logic_vector(31 downto 0);
    signal iNsTr_52_592 : std_logic_vector(31 downto 0);
    signal iNsTr_55_622 : std_logic_vector(31 downto 0);
    signal iNsTr_57_634 : std_logic_vector(31 downto 0);
    signal iNsTr_58_650 : std_logic_vector(31 downto 0);
    signal iNsTr_59_666 : std_logic_vector(31 downto 0);
    signal iNsTr_60_692 : std_logic_vector(31 downto 0);
    signal iNsTr_61_708 : std_logic_vector(31 downto 0);
    signal iNsTr_62_724 : std_logic_vector(31 downto 0);
    signal iNsTr_63_740 : std_logic_vector(31 downto 0);
    signal iNsTr_66_813 : std_logic_vector(63 downto 0);
    signal iNsTr_79_1020 : std_logic_vector(63 downto 0);
    signal iNsTr_81_1215 : std_logic_vector(31 downto 0);
    signal iNsTr_82_1231 : std_logic_vector(31 downto 0);
    signal iNsTr_83_1247 : std_logic_vector(31 downto 0);
    signal iNsTr_8_221 : std_logic_vector(31 downto 0);
    signal iNsTr_96_1300 : std_logic_vector(63 downto 0);
    signal inc63_286 : std_logic_vector(31 downto 0);
    signal inc_126 : std_logic_vector(31 downto 0);
    signal indvar332_1036 : std_logic_vector(63 downto 0);
    signal indvar348_829 : std_logic_vector(63 downto 0);
    signal indvar364_372 : std_logic_vector(63 downto 0);
    signal indvar367_269 : std_logic_vector(63 downto 0);
    signal indvar372_103 : std_logic_vector(63 downto 0);
    signal indvar_1316 : std_logic_vector(63 downto 0);
    signal indvarx_xnext333_1193 : std_logic_vector(63 downto 0);
    signal indvarx_xnext349_986 : std_logic_vector(63 downto 0);
    signal indvarx_xnext365_429 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1341 : std_logic_vector(63 downto 0);
    signal mul135_684 : std_logic_vector(31 downto 0);
    signal mul141_753 : std_logic_vector(31 downto 0);
    signal mul144_758 : std_logic_vector(31 downto 0);
    signal mul147_763 : std_logic_vector(31 downto 0);
    signal mul273_1260 : std_logic_vector(31 downto 0);
    signal mul276_1265 : std_logic_vector(31 downto 0);
    signal mul_679 : std_logic_vector(31 downto 0);
    signal ptr_deref_1185_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1185_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1185_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1185_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1185_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1185_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1218_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1218_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1218_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1218_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1218_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1234_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1234_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1234_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1234_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1234_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1250_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1250_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1250_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1250_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1250_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1332_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1332_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1332_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1332_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1332_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1332_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_135_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_135_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_135_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_135_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_135_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_135_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_157_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_157_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_157_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_157_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_157_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_157_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_174_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_174_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_174_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_174_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_174_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_223_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_223_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_223_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_223_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_223_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_223_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_251_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_251_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_251_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_251_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_251_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_251_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_302_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_302_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_302_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_302_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_302_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_302_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_324_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_324_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_324_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_324_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_324_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_324_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_341_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_341_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_341_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_341_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_341_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_392_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_392_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_392_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_392_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_392_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_392_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_414_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_414_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_414_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_414_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_414_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_414_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_496_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_496_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_496_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_496_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_496_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_496_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_49_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_49_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_49_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_49_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_49_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_49_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_526_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_526_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_526_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_526_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_526_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_526_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_545_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_545_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_545_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_545_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_545_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_545_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_575_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_575_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_575_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_575_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_575_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_575_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_594_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_594_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_594_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_594_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_594_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_594_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_624_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_624_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_624_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_624_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_624_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_624_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_637_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_637_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_637_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_637_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_637_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_653_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_653_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_653_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_653_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_653_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_669_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_669_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_669_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_669_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_669_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_695_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_695_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_695_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_695_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_695_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_711_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_711_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_711_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_711_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_711_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_727_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_727_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_727_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_727_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_727_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_743_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_743_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_743_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_743_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_743_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_77_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_77_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_77_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_77_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_77_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_77_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_978_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_978_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_978_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_978_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_978_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_978_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl105_504 : std_logic_vector(15 downto 0);
    signal shl114_553 : std_logic_vector(15 downto 0);
    signal shl123_602 : std_logic_vector(15 downto 0);
    signal shl158_856 : std_logic_vector(63 downto 0);
    signal shl164_874 : std_logic_vector(63 downto 0);
    signal shl170_892 : std_logic_vector(63 downto 0);
    signal shl176_910 : std_logic_vector(63 downto 0);
    signal shl182_928 : std_logic_vector(63 downto 0);
    signal shl188_946 : std_logic_vector(63 downto 0);
    signal shl18_143 : std_logic_vector(15 downto 0);
    signal shl194_964 : std_logic_vector(63 downto 0);
    signal shl219_1063 : std_logic_vector(63 downto 0);
    signal shl225_1081 : std_logic_vector(63 downto 0);
    signal shl231_1099 : std_logic_vector(63 downto 0);
    signal shl237_1117 : std_logic_vector(63 downto 0);
    signal shl243_1135 : std_logic_vector(63 downto 0);
    signal shl249_1153 : std_logic_vector(63 downto 0);
    signal shl255_1171 : std_logic_vector(63 downto 0);
    signal shl31_231 : std_logic_vector(15 downto 0);
    signal shl53_310 : std_logic_vector(15 downto 0);
    signal shl80_400 : std_logic_vector(15 downto 0);
    signal shl96_464 : std_logic_vector(15 downto 0);
    signal shl_57 : std_logic_vector(15 downto 0);
    signal tmp129_638 : std_logic_vector(15 downto 0);
    signal tmp131_654 : std_logic_vector(15 downto 0);
    signal tmp133_670 : std_logic_vector(15 downto 0);
    signal tmp137_696 : std_logic_vector(15 downto 0);
    signal tmp139_712 : std_logic_vector(15 downto 0);
    signal tmp142_728 : std_logic_vector(15 downto 0);
    signal tmp145_744 : std_logic_vector(15 downto 0);
    signal tmp269_1219 : std_logic_vector(15 downto 0);
    signal tmp271_1235 : std_logic_vector(15 downto 0);
    signal tmp274_1251 : std_logic_vector(15 downto 0);
    signal tmp327_1284 : std_logic_vector(31 downto 0);
    signal tmp327x_xop_1296 : std_logic_vector(31 downto 0);
    signal tmp328_1290 : std_logic_vector(0 downto 0);
    signal tmp331_1313 : std_logic_vector(63 downto 0);
    signal tmp341_1004 : std_logic_vector(31 downto 0);
    signal tmp341x_xop_1016 : std_logic_vector(31 downto 0);
    signal tmp342_1010 : std_logic_vector(0 downto 0);
    signal tmp346_1033 : std_logic_vector(63 downto 0);
    signal tmp355_797 : std_logic_vector(31 downto 0);
    signal tmp355x_xop_809 : std_logic_vector(31 downto 0);
    signal tmp356_803 : std_logic_vector(0 downto 0);
    signal tmp360_826 : std_logic_vector(63 downto 0);
    signal tmp369_332 : std_logic_vector(63 downto 0);
    signal tmp374_165 : std_logic_vector(63 downto 0);
    signal tmp38_342 : std_logic_vector(15 downto 0);
    signal tmp3_282 : std_logic_vector(63 downto 0);
    signal tmp7_175 : std_logic_vector(15 downto 0);
    signal tmp_122 : std_logic_vector(63 downto 0);
    signal type_cast_1002_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1008_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1014_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1024_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1031_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1040_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1042_wire : std_logic_vector(63 downto 0);
    signal type_cast_1061_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_106_wire : std_logic_vector(63 downto 0);
    signal type_cast_1079_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1097_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_109_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1115_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1133_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_113_wire : std_logic_vector(15 downto 0);
    signal type_cast_1151_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_115_wire : std_logic_vector(15 downto 0);
    signal type_cast_1169_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1191_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_120_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1269_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1282_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1288_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1294_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1304_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1311_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1320_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1322_wire : std_logic_vector(63 downto 0);
    signal type_cast_1334_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1339_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_141_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_163_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_183_wire : std_logic_vector(31 downto 0);
    signal type_cast_185_wire : std_logic_vector(31 downto 0);
    signal type_cast_205_wire : std_logic_vector(15 downto 0);
    signal type_cast_212_wire : std_logic_vector(15 downto 0);
    signal type_cast_214_wire : std_logic_vector(15 downto 0);
    signal type_cast_229_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_257_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_272_wire : std_logic_vector(63 downto 0);
    signal type_cast_275_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_280_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_308_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_330_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_349_wire : std_logic_vector(31 downto 0);
    signal type_cast_351_wire : std_logic_vector(31 downto 0);
    signal type_cast_376_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_378_wire : std_logic_vector(63 downto 0);
    signal type_cast_382_wire : std_logic_vector(15 downto 0);
    signal type_cast_384_wire : std_logic_vector(15 downto 0);
    signal type_cast_398_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_427_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_433_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_446_wire : std_logic_vector(15 downto 0);
    signal type_cast_450_wire : std_logic_vector(7 downto 0);
    signal type_cast_462_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_502_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_551_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_55_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_600_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_767_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_782_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_795_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_801_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_807_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_817_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_824_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_833_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_835_wire : std_logic_vector(63 downto 0);
    signal type_cast_83_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_854_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_872_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_890_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_908_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_926_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_944_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_962_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_984_wire_constant : std_logic_vector(63 downto 0);
    signal xx_xop376_1026 : std_logic_vector(63 downto 0);
    signal xx_xop377_819 : std_logic_vector(63 downto 0);
    signal xx_xop_1306 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_padding_452_word_address_0 <= "0";
    STORE_padding_477_word_address_0 <= "0";
    array_obj_ref_1048_constant_part_of_offset <= "00000010001";
    array_obj_ref_1048_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_1048_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_1048_resized_base_address <= "00000000000";
    array_obj_ref_131_constant_part_of_offset <= "0000100";
    array_obj_ref_131_offset_scale_factor_0 <= "1000000";
    array_obj_ref_131_offset_scale_factor_1 <= "0000001";
    array_obj_ref_131_resized_base_address <= "0000000";
    array_obj_ref_1328_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1328_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1328_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1328_resized_base_address <= "00000000000000";
    array_obj_ref_291_constant_part_of_offset <= "0000100";
    array_obj_ref_291_offset_scale_factor_0 <= "1000000";
    array_obj_ref_291_offset_scale_factor_1 <= "0000001";
    array_obj_ref_291_resized_base_address <= "0000000";
    array_obj_ref_388_offset_scale_factor_0 <= "1";
    array_obj_ref_388_resized_base_address <= "0";
    array_obj_ref_841_constant_part_of_offset <= "00000000000000";
    array_obj_ref_841_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_841_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_841_resized_base_address <= "00000000000000";
    iNsTr_11_249 <= "00000000000000000000000000000011";
    iNsTr_1_47 <= "00000000000000000000000000000011";
    iNsTr_21_171 <= "00000000000000000000000000000011";
    iNsTr_33_338 <= "00000000000000000000000000000011";
    iNsTr_40_494 <= "00000000000000000000000000000100";
    iNsTr_43_524 <= "00000000000000000000000000000100";
    iNsTr_46_543 <= "00000000000000000000000000000101";
    iNsTr_49_573 <= "00000000000000000000000000000101";
    iNsTr_4_75 <= "00000000000000000000000000000011";
    iNsTr_52_592 <= "00000000000000000000000000000110";
    iNsTr_55_622 <= "00000000000000000000000000000110";
    iNsTr_57_634 <= "00000000000000000000000000000100";
    iNsTr_58_650 <= "00000000000000000000000000000101";
    iNsTr_59_666 <= "00000000000000000000000000000110";
    iNsTr_60_692 <= "00000000000000000000000000000100";
    iNsTr_61_708 <= "00000000000000000000000000000101";
    iNsTr_62_724 <= "00000000000000000000000000000110";
    iNsTr_63_740 <= "00000000000000000000000000000111";
    iNsTr_81_1215 <= "00000000000000000000000000000100";
    iNsTr_82_1231 <= "00000000000000000000000000000101";
    iNsTr_83_1247 <= "00000000000000000000000000000110";
    iNsTr_8_221 <= "00000000000000000000000000000011";
    ptr_deref_1185_word_offset_0 <= "00000000000";
    ptr_deref_1218_word_offset_0 <= "0000000";
    ptr_deref_1234_word_offset_0 <= "0000000";
    ptr_deref_1250_word_offset_0 <= "0000000";
    ptr_deref_1332_word_offset_0 <= "00000000000000";
    ptr_deref_135_word_offset_0 <= "0000000";
    ptr_deref_157_word_offset_0 <= "0000000";
    ptr_deref_174_word_offset_0 <= "0000000";
    ptr_deref_223_word_offset_0 <= "0000000";
    ptr_deref_251_word_offset_0 <= "0000000";
    ptr_deref_302_word_offset_0 <= "0000000";
    ptr_deref_324_word_offset_0 <= "0000000";
    ptr_deref_341_word_offset_0 <= "0000000";
    ptr_deref_392_word_offset_0 <= "0";
    ptr_deref_414_word_offset_0 <= "0";
    ptr_deref_496_word_offset_0 <= "0000000";
    ptr_deref_49_word_offset_0 <= "0000000";
    ptr_deref_526_word_offset_0 <= "0000000";
    ptr_deref_545_word_offset_0 <= "0000000";
    ptr_deref_575_word_offset_0 <= "0000000";
    ptr_deref_594_word_offset_0 <= "0000000";
    ptr_deref_624_word_offset_0 <= "0000000";
    ptr_deref_637_word_offset_0 <= "0000000";
    ptr_deref_653_word_offset_0 <= "0000000";
    ptr_deref_669_word_offset_0 <= "0000000";
    ptr_deref_695_word_offset_0 <= "0000000";
    ptr_deref_711_word_offset_0 <= "0000000";
    ptr_deref_727_word_offset_0 <= "0000000";
    ptr_deref_743_word_offset_0 <= "0000000";
    ptr_deref_77_word_offset_0 <= "0000000";
    ptr_deref_978_word_offset_0 <= "00000000000000";
    type_cast_1002_wire_constant <= "00000000000000000000000000000010";
    type_cast_1008_wire_constant <= "00000000000000000000000000000001";
    type_cast_1014_wire_constant <= "11111111111111111111111111111111";
    type_cast_1024_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1031_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1040_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1061_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1079_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1097_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_109_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1115_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1133_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1151_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1169_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1191_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_120_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1269_wire_constant <= "00000000000000000000000000000011";
    type_cast_1282_wire_constant <= "00000000000000000000000000000010";
    type_cast_1288_wire_constant <= "00000000000000000000000000000001";
    type_cast_1294_wire_constant <= "11111111111111111111111111111111";
    type_cast_1304_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1311_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1320_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1334_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1339_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_141_wire_constant <= "0000000000001000";
    type_cast_163_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_229_wire_constant <= "0000000000001000";
    type_cast_257_wire_constant <= "0000000000000000";
    type_cast_275_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_280_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_308_wire_constant <= "0000000000001000";
    type_cast_330_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_376_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_398_wire_constant <= "0000000000001000";
    type_cast_427_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_433_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_462_wire_constant <= "0000000000001000";
    type_cast_502_wire_constant <= "0000000000001000";
    type_cast_551_wire_constant <= "0000000000001000";
    type_cast_55_wire_constant <= "0000000000001000";
    type_cast_600_wire_constant <= "0000000000001000";
    type_cast_767_wire_constant <= "00000000000000000000000000000011";
    type_cast_782_wire_constant <= "00000000000000000000000000000011";
    type_cast_795_wire_constant <= "00000000000000000000000000000010";
    type_cast_801_wire_constant <= "00000000000000000000000000000001";
    type_cast_807_wire_constant <= "11111111111111111111111111111111";
    type_cast_817_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_824_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_833_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_83_wire_constant <= "0000000000000000";
    type_cast_854_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_872_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_890_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_908_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_926_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_944_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_962_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_984_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_103: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_106_wire & type_cast_109_wire_constant;
      req <= phi_stmt_103_req_0 & phi_stmt_103_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_103",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_103_ack_0,
          idata => idata,
          odata => indvar372_103,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_103
    phi_stmt_1036: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1040_wire_constant & type_cast_1042_wire;
      req <= phi_stmt_1036_req_0 & phi_stmt_1036_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1036",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1036_ack_0,
          idata => idata,
          odata => indvar332_1036,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1036
    phi_stmt_110: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_113_wire & type_cast_115_wire;
      req <= phi_stmt_110_req_0 & phi_stmt_110_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_110",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_110_ack_0,
          idata => idata,
          odata => conv11320_110,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_110
    phi_stmt_1316: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1320_wire_constant & type_cast_1322_wire;
      req <= phi_stmt_1316_req_0 & phi_stmt_1316_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1316",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1316_ack_0,
          idata => idata,
          odata => indvar_1316,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1316
    phi_stmt_202: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_205_wire;
      req(0) <= phi_stmt_202_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_202",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_202_ack_0,
          idata => idata,
          odata => conv11x_xlcssa1_202,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_202
    phi_stmt_209: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_212_wire & type_cast_214_wire;
      req <= phi_stmt_209_req_0 & phi_stmt_209_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_209",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_209_ack_0,
          idata => idata,
          odata => conv11x_xlcssa_209,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_209
    phi_stmt_269: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_272_wire & type_cast_275_wire_constant;
      req <= phi_stmt_269_req_0 & phi_stmt_269_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_269",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_269_ack_0,
          idata => idata,
          odata => indvar367_269,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_269
    phi_stmt_372: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_376_wire_constant & type_cast_378_wire;
      req <= phi_stmt_372_req_0 & phi_stmt_372_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_372",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_372_ack_0,
          idata => idata,
          odata => indvar364_372,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_372
    phi_stmt_379: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_382_wire & type_cast_384_wire;
      req <= phi_stmt_379_req_0 & phi_stmt_379_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_379",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_379_ack_0,
          idata => idata,
          odata => conv71306_379,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_379
    phi_stmt_443: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_446_wire;
      req(0) <= phi_stmt_443_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_443",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_443_ack_0,
          idata => idata,
          odata => conv71x_xlcssa_443,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_443
    phi_stmt_447: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_450_wire;
      req(0) <= phi_stmt_447_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_447",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_447_ack_0,
          idata => idata,
          odata => call70x_xlcssa_447,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_447
    phi_stmt_829: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_833_wire_constant & type_cast_835_wire;
      req <= phi_stmt_829_req_0 & phi_stmt_829_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_829",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_829_ack_0,
          idata => idata,
          odata => indvar348_829,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_829
    -- flow-through select operator MUX_1032_inst
    tmp346_1033 <= xx_xop376_1026 when (tmp342_1010(0) /=  '0') else type_cast_1031_wire_constant;
    -- flow-through select operator MUX_1312_inst
    tmp331_1313 <= xx_xop_1306 when (tmp328_1290(0) /=  '0') else type_cast_1311_wire_constant;
    -- flow-through select operator MUX_825_inst
    tmp360_826 <= xx_xop377_819 when (tmp356_803(0) /=  '0') else type_cast_824_wire_constant;
    addr_of_1049_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1049_final_reg_req_0;
      addr_of_1049_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1049_final_reg_req_1;
      addr_of_1049_final_reg_ack_1<= rack(0);
      addr_of_1049_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1049_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1048_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx263_1050,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1329_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1329_final_reg_req_0;
      addr_of_1329_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1329_final_reg_req_1;
      addr_of_1329_final_reg_ack_1<= rack(0);
      addr_of_1329_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1329_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1328_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx286_1330,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_132_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_132_final_reg_req_0;
      addr_of_132_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_132_final_reg_req_1;
      addr_of_132_final_reg_ack_1<= rack(0);
      addr_of_132_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_132_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 7,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_131_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx25_133,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_292_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_292_final_reg_req_0;
      addr_of_292_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_292_final_reg_req_1;
      addr_of_292_final_reg_ack_1<= rack(0);
      addr_of_292_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_292_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 7,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_291_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx60_293,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_389_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_389_final_reg_req_0;
      addr_of_389_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_389_final_reg_req_1;
      addr_of_389_final_reg_ack_1<= rack(0);
      addr_of_389_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_389_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_388_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_390,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_842_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_842_final_reg_req_0;
      addr_of_842_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_842_final_reg_req_1;
      addr_of_842_final_reg_ack_1<= rack(0);
      addr_of_842_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_842_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_841_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx202_843,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1019_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1019_inst_req_0;
      type_cast_1019_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1019_inst_req_1;
      type_cast_1019_inst_ack_1<= rack(0);
      type_cast_1019_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1019_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp341x_xop_1016,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_79_1020,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1042_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1042_inst_req_0;
      type_cast_1042_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1042_inst_req_1;
      type_cast_1042_inst_ack_1<= rack(0);
      type_cast_1042_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1042_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext333_1193,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1042_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1056_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1056_inst_req_0;
      type_cast_1056_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1056_inst_req_1;
      type_cast_1056_inst_ack_1<= rack(0);
      type_cast_1056_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1056_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call216_1053,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv217_1057,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1069_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1069_inst_req_0;
      type_cast_1069_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1069_inst_req_1;
      type_cast_1069_inst_ack_1<= rack(0);
      type_cast_1069_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1069_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call220_1066,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv222_1070,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_106_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_106_inst_req_0;
      type_cast_106_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_106_inst_req_1;
      type_cast_106_inst_ack_1<= rack(0);
      type_cast_106_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_106_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp374_165,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_106_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1087_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1087_inst_req_0;
      type_cast_1087_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1087_inst_req_1;
      type_cast_1087_inst_ack_1<= rack(0);
      type_cast_1087_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1087_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call226_1084,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv228_1088,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1105_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1105_inst_req_0;
      type_cast_1105_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1105_inst_req_1;
      type_cast_1105_inst_ack_1<= rack(0);
      type_cast_1105_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1105_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call232_1102,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv234_1106,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1123_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1123_inst_req_0;
      type_cast_1123_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1123_inst_req_1;
      type_cast_1123_inst_ack_1<= rack(0);
      type_cast_1123_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1123_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call238_1120,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv240_1124,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_113_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_113_inst_req_0;
      type_cast_113_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_113_inst_req_1;
      type_cast_113_inst_ack_1<= rack(0);
      type_cast_113_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_113_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv11318_93,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_113_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1141_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1141_inst_req_0;
      type_cast_1141_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1141_inst_req_1;
      type_cast_1141_inst_ack_1<= rack(0);
      type_cast_1141_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1141_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call244_1138,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv246_1142,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1159_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1159_inst_req_0;
      type_cast_1159_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1159_inst_req_1;
      type_cast_1159_inst_ack_1<= rack(0);
      type_cast_1159_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1159_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call250_1156,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv252_1160,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_115_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_115_inst_req_0;
      type_cast_115_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_115_inst_req_1;
      type_cast_115_inst_ack_1<= rack(0);
      type_cast_115_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_115_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv11_194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_115_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1177_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1177_inst_req_0;
      type_cast_1177_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1177_inst_req_1;
      type_cast_1177_inst_ack_1<= rack(0);
      type_cast_1177_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1177_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call256_1174,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv258_1178,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1222_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1222_inst_req_0;
      type_cast_1222_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1222_inst_req_1;
      type_cast_1222_inst_ack_1<= rack(0);
      type_cast_1222_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1222_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp269_1219,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv270_1223,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1238_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1238_inst_req_0;
      type_cast_1238_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1238_inst_req_1;
      type_cast_1238_inst_ack_1<= rack(0);
      type_cast_1238_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1238_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp271_1235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv272_1239,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1254_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1254_inst_req_0;
      type_cast_1254_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1254_inst_req_1;
      type_cast_1254_inst_ack_1<= rack(0);
      type_cast_1254_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1254_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp274_1251,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv275_1255,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_125_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_125_inst_req_0;
      type_cast_125_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_125_inst_req_1;
      type_cast_125_inst_ack_1<= rack(0);
      type_cast_125_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_125_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_122,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc_126,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1299_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1299_inst_req_0;
      type_cast_1299_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1299_inst_req_1;
      type_cast_1299_inst_ack_1<= rack(0);
      type_cast_1299_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1299_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp327x_xop_1296,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_96_1300,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1322_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1322_inst_req_0;
      type_cast_1322_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1322_inst_req_1;
      type_cast_1322_inst_ack_1<= rack(0);
      type_cast_1322_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1322_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1341,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1322_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_149_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_149_inst_req_0;
      type_cast_149_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_149_inst_req_1;
      type_cast_149_inst_ack_1<= rack(0);
      type_cast_149_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_149_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_146,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_150,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_178_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_178_inst_req_0;
      type_cast_178_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_178_inst_req_1;
      type_cast_178_inst_ack_1<= rack(0);
      type_cast_178_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_178_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp7_175,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_179,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_183_inst
    process(inc_126) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := inc_126(31 downto 0);
      type_cast_183_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_185_inst
    process(conv8_179) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv8_179(31 downto 0);
      type_cast_185_wire <= tmp_var; -- 
    end process;
    type_cast_193_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_193_inst_req_0;
      type_cast_193_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_193_inst_req_1;
      type_cast_193_inst_ack_1<= rack(0);
      type_cast_193_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_193_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_190,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_194,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_205_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_205_inst_req_0;
      type_cast_205_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_205_inst_req_1;
      type_cast_205_inst_ack_1<= rack(0);
      type_cast_205_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_205_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv11_194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_205_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_212_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_212_inst_req_0;
      type_cast_212_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_212_inst_req_1;
      type_cast_212_inst_ack_1<= rack(0);
      type_cast_212_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_212_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv11318_93,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_212_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_214_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_214_inst_req_0;
      type_cast_214_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_214_inst_req_1;
      type_cast_214_inst_ack_1<= rack(0);
      type_cast_214_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_214_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv11x_xlcssa1_202,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_214_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_237_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_237_inst_req_0;
      type_cast_237_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_237_inst_req_1;
      type_cast_237_inst_ack_1<= rack(0);
      type_cast_237_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_237_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_234,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv33_238,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_272_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_272_inst_req_0;
      type_cast_272_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_272_inst_req_1;
      type_cast_272_inst_ack_1<= rack(0);
      type_cast_272_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_272_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp369_332,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_272_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_285_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_285_inst_req_0;
      type_cast_285_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_285_inst_req_1;
      type_cast_285_inst_ack_1<= rack(0);
      type_cast_285_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_285_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3_282,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc63_286,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_299_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_299_inst_req_0;
      type_cast_299_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_299_inst_req_1;
      type_cast_299_inst_ack_1<= rack(0);
      type_cast_299_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_299_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call43_296,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_300,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_316_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_316_inst_req_0;
      type_cast_316_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_316_inst_req_1;
      type_cast_316_inst_ack_1<= rack(0);
      type_cast_316_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_316_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call54_313,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv55_317,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_345_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_345_inst_req_0;
      type_cast_345_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_345_inst_req_1;
      type_cast_345_inst_ack_1<= rack(0);
      type_cast_345_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_345_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp38_342,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_346,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_349_inst
    process(inc63_286) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := inc63_286(31 downto 0);
      type_cast_349_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_351_inst
    process(conv39_346) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv39_346(31 downto 0);
      type_cast_351_wire <= tmp_var; -- 
    end process;
    type_cast_368_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_368_inst_req_0;
      type_cast_368_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_368_inst_req_1;
      type_cast_368_inst_ack_1<= rack(0);
      type_cast_368_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_368_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call70303_365,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71304_369,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_378_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_378_inst_req_0;
      type_cast_378_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_378_inst_req_1;
      type_cast_378_inst_ack_1<= rack(0);
      type_cast_378_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_378_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext365_429,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_378_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_382_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_382_inst_req_0;
      type_cast_382_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_382_inst_req_1;
      type_cast_382_inst_ack_1<= rack(0);
      type_cast_382_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_382_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv71304_369,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_382_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_384_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_384_inst_req_0;
      type_cast_384_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_384_inst_req_1;
      type_cast_384_inst_ack_1<= rack(0);
      type_cast_384_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_384_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv71_423,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_384_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_406_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_406_inst_req_0;
      type_cast_406_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_406_inst_req_1;
      type_cast_406_inst_ack_1<= rack(0);
      type_cast_406_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_406_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call81_403,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_407,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_40_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_40_inst_req_0;
      type_cast_40_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_40_inst_req_1;
      type_cast_40_inst_ack_1<= rack(0);
      type_cast_40_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_40_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_37,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_41,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_422_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_422_inst_req_0;
      type_cast_422_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_422_inst_req_1;
      type_cast_422_inst_ack_1<= rack(0);
      type_cast_422_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_422_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call70_419,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_423,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_446_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_446_inst_req_0;
      type_cast_446_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_446_inst_req_1;
      type_cast_446_inst_ack_1<= rack(0);
      type_cast_446_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_446_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv71_423,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_446_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_450_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_450_inst_req_0;
      type_cast_450_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_450_inst_req_1;
      type_cast_450_inst_ack_1<= rack(0);
      type_cast_450_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_450_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call70_419,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_450_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_457_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_457_inst_req_0;
      type_cast_457_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_457_inst_req_1;
      type_cast_457_inst_ack_1<= rack(0);
      type_cast_457_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_457_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call70x_xlcssa_447,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_458,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_470_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_470_inst_req_0;
      type_cast_470_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_470_inst_req_1;
      type_cast_470_inst_ack_1<= rack(0);
      type_cast_470_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_470_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_467,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_471,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_485_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_485_inst_req_0;
      type_cast_485_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_485_inst_req_1;
      type_cast_485_inst_ack_1<= rack(0);
      type_cast_485_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_485_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_482,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv102_486,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_510_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_510_inst_req_0;
      type_cast_510_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_510_inst_req_1;
      type_cast_510_inst_ack_1<= rack(0);
      type_cast_510_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_510_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_507,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_511,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_534_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_534_inst_req_0;
      type_cast_534_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_534_inst_req_1;
      type_cast_534_inst_ack_1<= rack(0);
      type_cast_534_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_534_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call110_531,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv111_535,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_559_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_559_inst_req_0;
      type_cast_559_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_559_inst_req_1;
      type_cast_559_inst_ack_1<= rack(0);
      type_cast_559_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_559_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_556,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_560,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_583_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_583_inst_req_0;
      type_cast_583_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_583_inst_req_1;
      type_cast_583_inst_ack_1<= rack(0);
      type_cast_583_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_583_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call119_580,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv120_584,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_608_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_608_inst_req_0;
      type_cast_608_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_608_inst_req_1;
      type_cast_608_inst_ack_1<= rack(0);
      type_cast_608_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_608_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call124_605,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_609,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_63_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_63_inst_req_0;
      type_cast_63_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_63_inst_req_1;
      type_cast_63_inst_ack_1<= rack(0);
      type_cast_63_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_63_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_60,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_64,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_641_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_641_inst_req_0;
      type_cast_641_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_641_inst_req_1;
      type_cast_641_inst_ack_1<= rack(0);
      type_cast_641_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_641_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp129_638,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv130_642,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_657_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_657_inst_req_0;
      type_cast_657_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_657_inst_req_1;
      type_cast_657_inst_ack_1<= rack(0);
      type_cast_657_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_657_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp131_654,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv132_658,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_673_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_673_inst_req_0;
      type_cast_673_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_673_inst_req_1;
      type_cast_673_inst_ack_1<= rack(0);
      type_cast_673_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_673_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp133_670,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_674,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_699_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_699_inst_req_0;
      type_cast_699_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_699_inst_req_1;
      type_cast_699_inst_ack_1<= rack(0);
      type_cast_699_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_699_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp137_696,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv138_700,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_715_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_715_inst_req_0;
      type_cast_715_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_715_inst_req_1;
      type_cast_715_inst_ack_1<= rack(0);
      type_cast_715_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_715_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp139_712,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv140_716,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_731_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_731_inst_req_0;
      type_cast_731_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_731_inst_req_1;
      type_cast_731_inst_ack_1<= rack(0);
      type_cast_731_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_731_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp142_728,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv143_732,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_747_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_747_inst_req_0;
      type_cast_747_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_747_inst_req_1;
      type_cast_747_inst_ack_1<= rack(0);
      type_cast_747_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_747_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp145_744,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv146_748,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_812_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_812_inst_req_0;
      type_cast_812_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_812_inst_req_1;
      type_cast_812_inst_ack_1<= rack(0);
      type_cast_812_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_812_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp355x_xop_809,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_66_813,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_835_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_835_inst_req_0;
      type_cast_835_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_835_inst_req_1;
      type_cast_835_inst_ack_1<= rack(0);
      type_cast_835_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_835_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext349_986,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_835_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_849_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_849_inst_req_0;
      type_cast_849_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_849_inst_req_1;
      type_cast_849_inst_ack_1<= rack(0);
      type_cast_849_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_849_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call155_846,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv156_850,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_862_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_862_inst_req_0;
      type_cast_862_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_862_inst_req_1;
      type_cast_862_inst_ack_1<= rack(0);
      type_cast_862_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_862_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call159_859,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv161_863,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_880_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_880_inst_req_0;
      type_cast_880_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_880_inst_req_1;
      type_cast_880_inst_ack_1<= rack(0);
      type_cast_880_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_880_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call165_877,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv167_881,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_898_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_898_inst_req_0;
      type_cast_898_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_898_inst_req_1;
      type_cast_898_inst_ack_1<= rack(0);
      type_cast_898_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_898_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call171_895,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv173_899,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_916_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_916_inst_req_0;
      type_cast_916_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_916_inst_req_1;
      type_cast_916_inst_ack_1<= rack(0);
      type_cast_916_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_916_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call177_913,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv179_917,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_92_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_92_inst_req_0;
      type_cast_92_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_92_inst_req_1;
      type_cast_92_inst_ack_1<= rack(0);
      type_cast_92_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_92_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10317_89,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11318_93,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_934_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_934_inst_req_0;
      type_cast_934_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_934_inst_req_1;
      type_cast_934_inst_ack_1<= rack(0);
      type_cast_934_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_934_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call183_931,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv185_935,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_952_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_952_inst_req_0;
      type_cast_952_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_952_inst_req_1;
      type_cast_952_inst_ack_1<= rack(0);
      type_cast_952_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_952_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call189_949,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv191_953,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_970_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_970_inst_req_0;
      type_cast_970_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_970_inst_req_1;
      type_cast_970_inst_ack_1<= rack(0);
      type_cast_970_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_970_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call195_967,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv197_971,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence STORE_padding_452_gather_scatter
    process(conv71x_xlcssa_443) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv71x_xlcssa_443;
      ov(15 downto 0) := iv;
      STORE_padding_452_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence STORE_padding_477_gather_scatter
    process(add99_476) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add99_476;
      ov(15 downto 0) := iv;
      STORE_padding_477_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1048_index_1_rename
    process(R_indvar332_1047_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar332_1047_resized;
      ov(10 downto 0) := iv;
      R_indvar332_1047_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1048_index_1_resize
    process(indvar332_1036) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar332_1036;
      ov := iv(10 downto 0);
      R_indvar332_1047_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1048_root_address_inst
    process(array_obj_ref_1048_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1048_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_1048_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_131_index_1_rename
    process(R_indvar372_130_resized) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar372_130_resized;
      ov(6 downto 0) := iv;
      R_indvar372_130_scaled <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_131_index_1_resize
    process(indvar372_103) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar372_103;
      ov := iv(6 downto 0);
      R_indvar372_130_resized <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_131_root_address_inst
    process(array_obj_ref_131_final_offset) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_131_final_offset;
      ov(6 downto 0) := iv;
      array_obj_ref_131_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1328_index_1_rename
    process(R_indvar_1327_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1327_resized;
      ov(13 downto 0) := iv;
      R_indvar_1327_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1328_index_1_resize
    process(indvar_1316) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1316;
      ov := iv(13 downto 0);
      R_indvar_1327_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1328_root_address_inst
    process(array_obj_ref_1328_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1328_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1328_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_291_index_1_rename
    process(R_indvar367_290_resized) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar367_290_resized;
      ov(6 downto 0) := iv;
      R_indvar367_290_scaled <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_291_index_1_resize
    process(indvar367_269) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar367_269;
      ov := iv(6 downto 0);
      R_indvar367_290_resized <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_291_root_address_inst
    process(array_obj_ref_291_final_offset) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_291_final_offset;
      ov(6 downto 0) := iv;
      array_obj_ref_291_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_388_index_0_rename
    process(R_indvar364_387_resized) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar364_387_resized;
      ov(0 downto 0) := iv;
      R_indvar364_387_scaled <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_388_index_0_resize
    process(indvar364_372) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar364_372;
      ov := iv(0 downto 0);
      R_indvar364_387_resized <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_388_index_offset
    process(R_indvar364_387_scaled) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar364_387_scaled;
      ov(0 downto 0) := iv;
      array_obj_ref_388_final_offset <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_388_root_address_inst
    process(array_obj_ref_388_final_offset) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_388_final_offset;
      ov(0 downto 0) := iv;
      array_obj_ref_388_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_841_index_1_rename
    process(R_indvar348_840_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar348_840_resized;
      ov(13 downto 0) := iv;
      R_indvar348_840_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_841_index_1_resize
    process(indvar348_829) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar348_829;
      ov := iv(13 downto 0);
      R_indvar348_840_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_841_root_address_inst
    process(array_obj_ref_841_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_841_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_841_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1185_addr_0
    process(ptr_deref_1185_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1185_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_1185_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1185_base_resize
    process(arrayidx263_1050) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx263_1050;
      ov := iv(10 downto 0);
      ptr_deref_1185_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1185_gather_scatter
    process(add259_1183) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add259_1183;
      ov(63 downto 0) := iv;
      ptr_deref_1185_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1185_root_address_inst
    process(ptr_deref_1185_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1185_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_1185_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1218_addr_0
    process(ptr_deref_1218_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1218_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1218_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1218_base_resize
    process(iNsTr_81_1215) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_81_1215;
      ov := iv(6 downto 0);
      ptr_deref_1218_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1218_gather_scatter
    process(ptr_deref_1218_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1218_data_0;
      ov(15 downto 0) := iv;
      tmp269_1219 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1218_root_address_inst
    process(ptr_deref_1218_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1218_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1218_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1234_addr_0
    process(ptr_deref_1234_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1234_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1234_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1234_base_resize
    process(iNsTr_82_1231) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_82_1231;
      ov := iv(6 downto 0);
      ptr_deref_1234_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1234_gather_scatter
    process(ptr_deref_1234_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1234_data_0;
      ov(15 downto 0) := iv;
      tmp271_1235 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1234_root_address_inst
    process(ptr_deref_1234_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1234_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1234_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1250_addr_0
    process(ptr_deref_1250_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1250_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1250_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1250_base_resize
    process(iNsTr_83_1247) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_83_1247;
      ov := iv(6 downto 0);
      ptr_deref_1250_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1250_gather_scatter
    process(ptr_deref_1250_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1250_data_0;
      ov(15 downto 0) := iv;
      tmp274_1251 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1250_root_address_inst
    process(ptr_deref_1250_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1250_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1250_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1332_addr_0
    process(ptr_deref_1332_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1332_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1332_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1332_base_resize
    process(arrayidx286_1330) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx286_1330;
      ov := iv(13 downto 0);
      ptr_deref_1332_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1332_gather_scatter
    process(type_cast_1334_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1334_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1332_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1332_root_address_inst
    process(ptr_deref_1332_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1332_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1332_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_135_addr_0
    process(ptr_deref_135_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_135_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_135_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_135_base_resize
    process(arrayidx25_133) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx25_133;
      ov := iv(6 downto 0);
      ptr_deref_135_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_135_gather_scatter
    process(conv11320_110) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv11320_110;
      ov(15 downto 0) := iv;
      ptr_deref_135_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_135_root_address_inst
    process(ptr_deref_135_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_135_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_135_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_157_addr_0
    process(ptr_deref_157_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_157_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_157_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_157_base_resize
    process(arrayidx25_133) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx25_133;
      ov := iv(6 downto 0);
      ptr_deref_157_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_157_gather_scatter
    process(add21_155) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add21_155;
      ov(15 downto 0) := iv;
      ptr_deref_157_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_157_root_address_inst
    process(ptr_deref_157_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_157_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_157_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_174_addr_0
    process(ptr_deref_174_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_174_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_174_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_174_base_resize
    process(iNsTr_21_171) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_21_171;
      ov := iv(6 downto 0);
      ptr_deref_174_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_174_gather_scatter
    process(ptr_deref_174_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_174_data_0;
      ov(15 downto 0) := iv;
      tmp7_175 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_174_root_address_inst
    process(ptr_deref_174_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_174_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_174_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_223_addr_0
    process(ptr_deref_223_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_223_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_223_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_223_base_resize
    process(iNsTr_8_221) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_221;
      ov := iv(6 downto 0);
      ptr_deref_223_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_223_gather_scatter
    process(conv11x_xlcssa_209) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv11x_xlcssa_209;
      ov(15 downto 0) := iv;
      ptr_deref_223_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_223_root_address_inst
    process(ptr_deref_223_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_223_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_223_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_251_addr_0
    process(ptr_deref_251_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_251_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_251_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_251_base_resize
    process(iNsTr_11_249) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_11_249;
      ov := iv(6 downto 0);
      ptr_deref_251_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_251_gather_scatter
    process(add34_243) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add34_243;
      ov(15 downto 0) := iv;
      ptr_deref_251_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_251_root_address_inst
    process(ptr_deref_251_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_251_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_251_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_302_addr_0
    process(ptr_deref_302_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_302_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_302_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_302_base_resize
    process(arrayidx60_293) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx60_293;
      ov := iv(6 downto 0);
      ptr_deref_302_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_302_gather_scatter
    process(conv44_300) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv44_300;
      ov(15 downto 0) := iv;
      ptr_deref_302_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_302_root_address_inst
    process(ptr_deref_302_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_302_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_302_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_324_addr_0
    process(ptr_deref_324_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_324_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_324_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_324_base_resize
    process(arrayidx60_293) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx60_293;
      ov := iv(6 downto 0);
      ptr_deref_324_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_324_gather_scatter
    process(add56_322) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add56_322;
      ov(15 downto 0) := iv;
      ptr_deref_324_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_324_root_address_inst
    process(ptr_deref_324_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_324_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_324_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_341_addr_0
    process(ptr_deref_341_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_341_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_341_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_341_base_resize
    process(iNsTr_33_338) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_33_338;
      ov := iv(6 downto 0);
      ptr_deref_341_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_341_gather_scatter
    process(ptr_deref_341_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_341_data_0;
      ov(15 downto 0) := iv;
      tmp38_342 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_341_root_address_inst
    process(ptr_deref_341_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_341_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_341_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_392_addr_0
    process(ptr_deref_392_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_392_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_392_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_392_base_resize
    process(arrayidx87_390) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_390;
      ov := iv(0 downto 0);
      ptr_deref_392_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_392_gather_scatter
    process(conv71306_379) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv71306_379;
      ov(15 downto 0) := iv;
      ptr_deref_392_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_392_root_address_inst
    process(ptr_deref_392_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_392_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_392_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_414_addr_0
    process(ptr_deref_414_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_414_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_414_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_414_base_resize
    process(arrayidx87_390) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_390;
      ov := iv(0 downto 0);
      ptr_deref_414_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_414_gather_scatter
    process(add83_412) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add83_412;
      ov(15 downto 0) := iv;
      ptr_deref_414_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_414_root_address_inst
    process(ptr_deref_414_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_414_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_414_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_496_addr_0
    process(ptr_deref_496_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_496_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_496_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_496_base_resize
    process(iNsTr_40_494) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_40_494;
      ov := iv(6 downto 0);
      ptr_deref_496_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_496_gather_scatter
    process(conv102_486) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv102_486;
      ov(15 downto 0) := iv;
      ptr_deref_496_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_496_root_address_inst
    process(ptr_deref_496_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_496_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_496_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_49_addr_0
    process(ptr_deref_49_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_49_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_49_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_49_base_resize
    process(iNsTr_1_47) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_1_47;
      ov := iv(6 downto 0);
      ptr_deref_49_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_49_gather_scatter
    process(conv_41) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv_41;
      ov(15 downto 0) := iv;
      ptr_deref_49_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_49_root_address_inst
    process(ptr_deref_49_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_49_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_49_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_526_addr_0
    process(ptr_deref_526_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_526_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_526_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_526_base_resize
    process(iNsTr_43_524) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_43_524;
      ov := iv(6 downto 0);
      ptr_deref_526_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_526_gather_scatter
    process(add108_516) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add108_516;
      ov(15 downto 0) := iv;
      ptr_deref_526_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_526_root_address_inst
    process(ptr_deref_526_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_526_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_526_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_545_addr_0
    process(ptr_deref_545_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_545_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_545_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_545_base_resize
    process(iNsTr_46_543) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_46_543;
      ov := iv(6 downto 0);
      ptr_deref_545_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_545_gather_scatter
    process(conv111_535) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv111_535;
      ov(15 downto 0) := iv;
      ptr_deref_545_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_545_root_address_inst
    process(ptr_deref_545_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_545_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_545_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_575_addr_0
    process(ptr_deref_575_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_575_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_575_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_575_base_resize
    process(iNsTr_49_573) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_49_573;
      ov := iv(6 downto 0);
      ptr_deref_575_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_575_gather_scatter
    process(add117_565) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add117_565;
      ov(15 downto 0) := iv;
      ptr_deref_575_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_575_root_address_inst
    process(ptr_deref_575_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_575_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_575_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_594_addr_0
    process(ptr_deref_594_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_594_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_594_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_594_base_resize
    process(iNsTr_52_592) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_52_592;
      ov := iv(6 downto 0);
      ptr_deref_594_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_594_gather_scatter
    process(conv120_584) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv120_584;
      ov(15 downto 0) := iv;
      ptr_deref_594_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_594_root_address_inst
    process(ptr_deref_594_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_594_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_594_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_624_addr_0
    process(ptr_deref_624_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_624_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_624_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_624_base_resize
    process(iNsTr_55_622) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_55_622;
      ov := iv(6 downto 0);
      ptr_deref_624_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_624_gather_scatter
    process(add126_614) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add126_614;
      ov(15 downto 0) := iv;
      ptr_deref_624_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_624_root_address_inst
    process(ptr_deref_624_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_624_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_624_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_637_addr_0
    process(ptr_deref_637_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_637_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_637_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_637_base_resize
    process(iNsTr_57_634) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_57_634;
      ov := iv(6 downto 0);
      ptr_deref_637_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_637_gather_scatter
    process(ptr_deref_637_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_637_data_0;
      ov(15 downto 0) := iv;
      tmp129_638 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_637_root_address_inst
    process(ptr_deref_637_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_637_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_637_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_653_addr_0
    process(ptr_deref_653_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_653_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_653_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_653_base_resize
    process(iNsTr_58_650) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_58_650;
      ov := iv(6 downto 0);
      ptr_deref_653_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_653_gather_scatter
    process(ptr_deref_653_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_653_data_0;
      ov(15 downto 0) := iv;
      tmp131_654 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_653_root_address_inst
    process(ptr_deref_653_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_653_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_653_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_669_addr_0
    process(ptr_deref_669_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_669_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_669_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_669_base_resize
    process(iNsTr_59_666) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_59_666;
      ov := iv(6 downto 0);
      ptr_deref_669_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_669_gather_scatter
    process(ptr_deref_669_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_669_data_0;
      ov(15 downto 0) := iv;
      tmp133_670 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_669_root_address_inst
    process(ptr_deref_669_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_669_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_669_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_695_addr_0
    process(ptr_deref_695_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_695_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_695_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_695_base_resize
    process(iNsTr_60_692) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_60_692;
      ov := iv(6 downto 0);
      ptr_deref_695_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_695_gather_scatter
    process(ptr_deref_695_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_695_data_0;
      ov(15 downto 0) := iv;
      tmp137_696 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_695_root_address_inst
    process(ptr_deref_695_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_695_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_695_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_711_addr_0
    process(ptr_deref_711_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_711_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_711_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_711_base_resize
    process(iNsTr_61_708) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_61_708;
      ov := iv(6 downto 0);
      ptr_deref_711_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_711_gather_scatter
    process(ptr_deref_711_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_711_data_0;
      ov(15 downto 0) := iv;
      tmp139_712 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_711_root_address_inst
    process(ptr_deref_711_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_711_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_711_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_727_addr_0
    process(ptr_deref_727_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_727_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_727_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_727_base_resize
    process(iNsTr_62_724) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_62_724;
      ov := iv(6 downto 0);
      ptr_deref_727_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_727_gather_scatter
    process(ptr_deref_727_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_727_data_0;
      ov(15 downto 0) := iv;
      tmp142_728 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_727_root_address_inst
    process(ptr_deref_727_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_727_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_727_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_743_addr_0
    process(ptr_deref_743_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_743_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_743_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_743_base_resize
    process(iNsTr_63_740) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_63_740;
      ov := iv(6 downto 0);
      ptr_deref_743_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_743_gather_scatter
    process(ptr_deref_743_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_743_data_0;
      ov(15 downto 0) := iv;
      tmp145_744 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_743_root_address_inst
    process(ptr_deref_743_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_743_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_743_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_77_addr_0
    process(ptr_deref_77_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_77_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_77_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_77_base_resize
    process(iNsTr_4_75) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_75;
      ov := iv(6 downto 0);
      ptr_deref_77_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_77_gather_scatter
    process(add_69) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add_69;
      ov(15 downto 0) := iv;
      ptr_deref_77_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_77_root_address_inst
    process(ptr_deref_77_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_77_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_77_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_978_addr_0
    process(ptr_deref_978_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_978_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_978_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_978_base_resize
    process(arrayidx202_843) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx202_843;
      ov := iv(13 downto 0);
      ptr_deref_978_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_978_gather_scatter
    process(add198_976) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add198_976;
      ov(63 downto 0) := iv;
      ptr_deref_978_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_978_root_address_inst
    process(ptr_deref_978_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_978_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_978_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1199_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_1198;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1199_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1199_branch_req_0,
          ack0 => if_stmt_1199_branch_ack_0,
          ack1 => if_stmt_1199_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1272_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp281292_1271;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1272_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1272_branch_req_0,
          ack0 => if_stmt_1272_branch_ack_0,
          ack1 => if_stmt_1272_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1347_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond5_1346;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1347_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1347_branch_req_0,
          ack0 => if_stmt_1347_branch_ack_0,
          ack1 => if_stmt_1347_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_195_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_187;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_195_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_195_branch_req_0,
          ack0 => if_stmt_195_branch_ack_0,
          ack1 => if_stmt_195_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_260_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp40311_259;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_260_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_260_branch_req_0,
          ack0 => if_stmt_260_branch_ack_0,
          ack1 => if_stmt_260_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_354_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp40_353;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_354_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_354_branch_req_0,
          ack0 => if_stmt_354_branch_ack_0,
          ack1 => if_stmt_354_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_436_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond7_435;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_436_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_436_branch_req_0,
          ack0 => if_stmt_436_branch_ack_0,
          ack1 => if_stmt_436_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_770_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp151299_769;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_770_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_770_branch_req_0,
          ack0 => if_stmt_770_branch_ack_0,
          ack1 => if_stmt_770_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_785_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp211295_784;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_785_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_785_branch_req_0,
          ack0 => if_stmt_785_branch_ack_0,
          ack1 => if_stmt_785_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_94_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp316_86;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_94_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_94_branch_req_0,
          ack0 => if_stmt_94_branch_ack_0,
          ack1 => if_stmt_94_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_992_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond6_991;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_992_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_992_branch_req_0,
          ack0 => if_stmt_992_branch_ack_0,
          ack1 => if_stmt_992_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1015_inst
    process(tmp341_1004) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp341_1004, type_cast_1014_wire_constant, tmp_var);
      tmp341x_xop_1016 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1295_inst
    process(tmp327_1284) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp327_1284, type_cast_1294_wire_constant, tmp_var);
      tmp327x_xop_1296 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_808_inst
    process(tmp355_797) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp355_797, type_cast_807_wire_constant, tmp_var);
      tmp355x_xop_809 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1025_inst
    process(iNsTr_79_1020) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_79_1020, type_cast_1024_wire_constant, tmp_var);
      xx_xop376_1026 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1192_inst
    process(indvar332_1036) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar332_1036, type_cast_1191_wire_constant, tmp_var);
      indvarx_xnext333_1193 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_121_inst
    process(indvar372_103) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar372_103, type_cast_120_wire_constant, tmp_var);
      tmp_122 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1305_inst
    process(iNsTr_96_1300) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_96_1300, type_cast_1304_wire_constant, tmp_var);
      xx_xop_1306 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1340_inst
    process(indvar_1316) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1316, type_cast_1339_wire_constant, tmp_var);
      indvarx_xnext_1341 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_164_inst
    process(indvar372_103) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar372_103, type_cast_163_wire_constant, tmp_var);
      tmp374_165 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_281_inst
    process(indvar367_269) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar367_269, type_cast_280_wire_constant, tmp_var);
      tmp3_282 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_331_inst
    process(indvar367_269) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar367_269, type_cast_330_wire_constant, tmp_var);
      tmp369_332 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_428_inst
    process(indvar364_372) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar364_372, type_cast_427_wire_constant, tmp_var);
      indvarx_xnext365_429 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_818_inst
    process(iNsTr_66_813) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_66_813, type_cast_817_wire_constant, tmp_var);
      xx_xop377_819 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_985_inst
    process(indvar348_829) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar348_829, type_cast_984_wire_constant, tmp_var);
      indvarx_xnext349_986 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_258_inst
    process(add34_243) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(add34_243, type_cast_257_wire_constant, tmp_var);
      cmp40311_259 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_84_inst
    process(add_69) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(add_69, type_cast_83_wire_constant, tmp_var);
      cmp316_86 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1197_inst
    process(indvarx_xnext333_1193, tmp346_1033) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext333_1193, tmp346_1033, tmp_var);
      exitcond_1198 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1345_inst
    process(indvarx_xnext_1341, tmp331_1313) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1341, tmp331_1313, tmp_var);
      exitcond5_1346 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_434_inst
    process(indvarx_xnext365_429) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext365_429, type_cast_433_wire_constant, tmp_var);
      exitcond7_435 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_990_inst
    process(indvarx_xnext349_986, tmp360_826) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext349_986, tmp360_826, tmp_var);
      exitcond6_991 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1003_inst
    process(mul147_763) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul147_763, type_cast_1002_wire_constant, tmp_var);
      tmp341_1004 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1283_inst
    process(mul276_1265) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul276_1265, type_cast_1282_wire_constant, tmp_var);
      tmp327_1284 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_796_inst
    process(mul135_684) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul135_684, type_cast_795_wire_constant, tmp_var);
      tmp355_797 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1259_inst
    process(conv272_1239, conv270_1223) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv272_1239, conv270_1223, tmp_var);
      mul273_1260 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1264_inst
    process(mul273_1260, conv275_1255) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul273_1260, conv275_1255, tmp_var);
      mul276_1265 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_678_inst
    process(conv132_658, conv130_642) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv132_658, conv130_642, tmp_var);
      mul_679 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_683_inst
    process(mul_679, conv134_674) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_679, conv134_674, tmp_var);
      mul135_684 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_752_inst
    process(conv140_716, conv138_700) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv140_716, conv138_700, tmp_var);
      mul141_753 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_757_inst
    process(mul141_753, conv143_732) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul141_753, conv143_732, tmp_var);
      mul144_758 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_762_inst
    process(mul144_758, conv146_748) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul144_758, conv146_748, tmp_var);
      mul147_763 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_154_inst
    process(conv20_150, shl18_143) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv20_150, shl18_143, tmp_var);
      add21_155 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_242_inst
    process(conv33_238, shl31_231) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv33_238, shl31_231, tmp_var);
      add34_243 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_321_inst
    process(conv55_317, shl53_310) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv55_317, shl53_310, tmp_var);
      add56_322 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_411_inst
    process(conv82_407, shl80_400) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv82_407, shl80_400, tmp_var);
      add83_412 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_475_inst
    process(conv98_471, shl96_464) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv98_471, shl96_464, tmp_var);
      add99_476 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_515_inst
    process(shl105_504, conv107_511) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl105_504, conv107_511, tmp_var);
      add108_516 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_564_inst
    process(shl114_553, conv116_560) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl114_553, conv116_560, tmp_var);
      add117_565 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_613_inst
    process(shl123_602, conv125_609) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl123_602, conv125_609, tmp_var);
      add126_614 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_68_inst
    process(shl_57, conv3_64) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_57, conv3_64, tmp_var);
      add_69 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1074_inst
    process(shl219_1063, conv222_1070) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl219_1063, conv222_1070, tmp_var);
      add223_1075 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1092_inst
    process(shl225_1081, conv228_1088) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl225_1081, conv228_1088, tmp_var);
      add229_1093 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1110_inst
    process(shl231_1099, conv234_1106) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl231_1099, conv234_1106, tmp_var);
      add235_1111 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1128_inst
    process(shl237_1117, conv240_1124) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl237_1117, conv240_1124, tmp_var);
      add241_1129 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1146_inst
    process(shl243_1135, conv246_1142) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl243_1135, conv246_1142, tmp_var);
      add247_1147 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1164_inst
    process(shl249_1153, conv252_1160) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl249_1153, conv252_1160, tmp_var);
      add253_1165 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1182_inst
    process(shl255_1171, conv258_1178) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl255_1171, conv258_1178, tmp_var);
      add259_1183 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_867_inst
    process(shl158_856, conv161_863) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl158_856, conv161_863, tmp_var);
      add162_868 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_885_inst
    process(shl164_874, conv167_881) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl164_874, conv167_881, tmp_var);
      add168_886 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_903_inst
    process(shl170_892, conv173_899) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl170_892, conv173_899, tmp_var);
      add174_904 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_921_inst
    process(shl176_910, conv179_917) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl176_910, conv179_917, tmp_var);
      add180_922 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_939_inst
    process(shl182_928, conv185_935) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl182_928, conv185_935, tmp_var);
      add186_940 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_957_inst
    process(shl188_946, conv191_953) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl188_946, conv191_953, tmp_var);
      add192_958 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_975_inst
    process(shl194_964, conv197_971) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl194_964, conv197_971, tmp_var);
      add198_976 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_142_inst
    process(conv11320_110) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv11320_110, type_cast_141_wire_constant, tmp_var);
      shl18_143 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_230_inst
    process(conv11x_xlcssa_209) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv11x_xlcssa_209, type_cast_229_wire_constant, tmp_var);
      shl31_231 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_309_inst
    process(conv44_300) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_300, type_cast_308_wire_constant, tmp_var);
      shl53_310 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_399_inst
    process(conv71306_379) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv71306_379, type_cast_398_wire_constant, tmp_var);
      shl80_400 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_463_inst
    process(conv95_458) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv95_458, type_cast_462_wire_constant, tmp_var);
      shl96_464 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_503_inst
    process(conv102_486) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv102_486, type_cast_502_wire_constant, tmp_var);
      shl105_504 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_552_inst
    process(conv111_535) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv111_535, type_cast_551_wire_constant, tmp_var);
      shl114_553 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_56_inst
    process(conv_41) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_41, type_cast_55_wire_constant, tmp_var);
      shl_57 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_601_inst
    process(conv120_584) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv120_584, type_cast_600_wire_constant, tmp_var);
      shl123_602 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1062_inst
    process(conv217_1057) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv217_1057, type_cast_1061_wire_constant, tmp_var);
      shl219_1063 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1080_inst
    process(add223_1075) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add223_1075, type_cast_1079_wire_constant, tmp_var);
      shl225_1081 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1098_inst
    process(add229_1093) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add229_1093, type_cast_1097_wire_constant, tmp_var);
      shl231_1099 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1116_inst
    process(add235_1111) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add235_1111, type_cast_1115_wire_constant, tmp_var);
      shl237_1117 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1134_inst
    process(add241_1129) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add241_1129, type_cast_1133_wire_constant, tmp_var);
      shl243_1135 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1152_inst
    process(add247_1147) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add247_1147, type_cast_1151_wire_constant, tmp_var);
      shl249_1153 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1170_inst
    process(add253_1165) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add253_1165, type_cast_1169_wire_constant, tmp_var);
      shl255_1171 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_855_inst
    process(conv156_850) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv156_850, type_cast_854_wire_constant, tmp_var);
      shl158_856 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_873_inst
    process(add162_868) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add162_868, type_cast_872_wire_constant, tmp_var);
      shl164_874 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_891_inst
    process(add168_886) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add168_886, type_cast_890_wire_constant, tmp_var);
      shl170_892 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_909_inst
    process(add174_904) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add174_904, type_cast_908_wire_constant, tmp_var);
      shl176_910 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_927_inst
    process(add180_922) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add180_922, type_cast_926_wire_constant, tmp_var);
      shl182_928 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_945_inst
    process(add186_940) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add186_940, type_cast_944_wire_constant, tmp_var);
      shl188_946 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_963_inst
    process(add192_958) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add192_958, type_cast_962_wire_constant, tmp_var);
      shl194_964 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_186_inst
    process(type_cast_183_wire, type_cast_185_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_183_wire, type_cast_185_wire, tmp_var);
      cmp_187 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_352_inst
    process(type_cast_349_wire, type_cast_351_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_349_wire, type_cast_351_wire, tmp_var);
      cmp40_353 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1009_inst
    process(tmp341_1004) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp341_1004, type_cast_1008_wire_constant, tmp_var);
      tmp342_1010 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1270_inst
    process(mul276_1265) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul276_1265, type_cast_1269_wire_constant, tmp_var);
      cmp281292_1271 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1289_inst
    process(tmp327_1284) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp327_1284, type_cast_1288_wire_constant, tmp_var);
      tmp328_1290 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_768_inst
    process(mul135_684) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul135_684, type_cast_767_wire_constant, tmp_var);
      cmp151299_769 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_783_inst
    process(mul147_763) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul147_763, type_cast_782_wire_constant, tmp_var);
      cmp211295_784 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_802_inst
    process(tmp355_797) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp355_797, type_cast_801_wire_constant, tmp_var);
      tmp356_803 <= tmp_var; --
    end process;
    -- shared split operator group (84) : array_obj_ref_1048_index_offset 
    ApIntAdd_group_84: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar332_1047_scaled;
      array_obj_ref_1048_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1048_index_offset_req_0;
      array_obj_ref_1048_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1048_index_offset_req_1;
      array_obj_ref_1048_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_84_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_84_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_84",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000010001",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 84
    -- shared split operator group (85) : array_obj_ref_131_index_offset 
    ApIntAdd_group_85: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(6 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar372_130_scaled;
      array_obj_ref_131_final_offset <= data_out(6 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_131_index_offset_req_0;
      array_obj_ref_131_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_131_index_offset_req_1;
      array_obj_ref_131_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_85_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_85_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_85",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0000100",
          constant_width => 7,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 85
    -- shared split operator group (86) : array_obj_ref_1328_index_offset 
    ApIntAdd_group_86: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1327_scaled;
      array_obj_ref_1328_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1328_index_offset_req_0;
      array_obj_ref_1328_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1328_index_offset_req_1;
      array_obj_ref_1328_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_86_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_86_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_86",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 86
    -- shared split operator group (87) : array_obj_ref_291_index_offset 
    ApIntAdd_group_87: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(6 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar367_290_scaled;
      array_obj_ref_291_final_offset <= data_out(6 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_291_index_offset_req_0;
      array_obj_ref_291_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_291_index_offset_req_1;
      array_obj_ref_291_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_87_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_87_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_87",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0000100",
          constant_width => 7,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 87
    -- shared split operator group (88) : array_obj_ref_841_index_offset 
    ApIntAdd_group_88: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar348_840_scaled;
      array_obj_ref_841_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_841_index_offset_req_0;
      array_obj_ref_841_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_841_index_offset_req_1;
      array_obj_ref_841_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_88_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_88_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_88",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 88
    -- shared load operator group (0) : ptr_deref_1218_load_0 ptr_deref_1234_load_0 ptr_deref_1250_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1218_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1234_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1250_load_0_req_0;
      ptr_deref_1218_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1234_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1250_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1218_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1234_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1250_load_0_req_1;
      ptr_deref_1218_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1234_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1250_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1218_word_address_0 & ptr_deref_1234_word_address_0 & ptr_deref_1250_word_address_0;
      ptr_deref_1218_data_0 <= data_out(47 downto 32);
      ptr_deref_1234_data_0 <= data_out(31 downto 16);
      ptr_deref_1250_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(15 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_669_load_0 ptr_deref_653_load_0 ptr_deref_637_load_0 ptr_deref_174_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_669_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_653_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_637_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_174_load_0_req_0;
      ptr_deref_669_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_653_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_637_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_174_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_669_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_653_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_637_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_174_load_0_req_1;
      ptr_deref_669_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_653_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_637_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_174_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_669_word_address_0 & ptr_deref_653_word_address_0 & ptr_deref_637_word_address_0 & ptr_deref_174_word_address_0;
      ptr_deref_669_data_0 <= data_out(63 downto 48);
      ptr_deref_653_data_0 <= data_out(47 downto 32);
      ptr_deref_637_data_0 <= data_out(31 downto 16);
      ptr_deref_174_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 16,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(15 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_341_load_0 ptr_deref_695_load_0 ptr_deref_711_load_0 ptr_deref_727_load_0 ptr_deref_743_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(34 downto 0);
      signal data_out: std_logic_vector(79 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 4 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 4 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 4 downto 0);
      signal guard_vector : std_logic_vector( 4 downto 0);
      constant inBUFs : IntegerArray(4 downto 0) := (4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(4 downto 0) := (4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(4 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false);
      constant guardBuffering: IntegerArray(4 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2);
      -- 
    begin -- 
      reqL_unguarded(4) <= ptr_deref_341_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_695_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_711_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_727_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_743_load_0_req_0;
      ptr_deref_341_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_695_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_711_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_727_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_743_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(4) <= ptr_deref_341_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_695_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_711_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_727_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_743_load_0_req_1;
      ptr_deref_341_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_695_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_711_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_727_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_743_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 5, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_341_word_address_0 & ptr_deref_695_word_address_0 & ptr_deref_711_word_address_0 & ptr_deref_727_word_address_0 & ptr_deref_743_word_address_0;
      ptr_deref_341_data_0 <= data_out(79 downto 64);
      ptr_deref_695_data_0 <= data_out(63 downto 48);
      ptr_deref_711_data_0 <= data_out(47 downto 32);
      ptr_deref_727_data_0 <= data_out(31 downto 16);
      ptr_deref_743_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 7,
        num_reqs => 5,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 5,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(15 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared store operator group (0) : STORE_padding_477_store_0 STORE_padding_452_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(1 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= STORE_padding_477_store_0_req_0;
      reqL_unguarded(0) <= STORE_padding_452_store_0_req_0;
      STORE_padding_477_store_0_ack_0 <= ackL_unguarded(1);
      STORE_padding_452_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= STORE_padding_477_store_0_req_1;
      reqR_unguarded(0) <= STORE_padding_452_store_0_req_1;
      STORE_padding_477_store_0_ack_1 <= ackR_unguarded(1);
      STORE_padding_452_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_padding_477_word_address_0 & STORE_padding_452_word_address_0;
      data_in <= STORE_padding_477_data_0 & STORE_padding_452_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_7_sr_req(0),
          mack => memory_space_7_sr_ack(0),
          maddr => memory_space_7_sr_addr(0 downto 0),
          mdata => memory_space_7_sr_data(15 downto 0),
          mtag => memory_space_7_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_7_sc_req(0),
          mack => memory_space_7_sc_ack(0),
          mtag => memory_space_7_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_1185_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1185_store_0_req_0;
      ptr_deref_1185_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1185_store_0_req_1;
      ptr_deref_1185_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1185_word_address_0;
      data_in <= ptr_deref_1185_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(10 downto 0),
          mdata => memory_space_5_sr_data(63 downto 0),
          mtag => memory_space_5_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_1332_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1332_store_0_req_0;
      ptr_deref_1332_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1332_store_0_req_1;
      ptr_deref_1332_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1332_word_address_0;
      data_in <= ptr_deref_1332_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(13 downto 0),
          mdata => memory_space_6_sr_data(63 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_49_store_0 ptr_deref_77_store_0 ptr_deref_135_store_0 ptr_deref_157_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_49_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_77_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_135_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_157_store_0_req_0;
      ptr_deref_49_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_77_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_135_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_157_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_49_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_77_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_135_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_157_store_0_req_1;
      ptr_deref_49_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_77_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_135_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_157_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      StoreGroup3_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_49_word_address_0 & ptr_deref_77_word_address_0 & ptr_deref_135_word_address_0 & ptr_deref_157_word_address_0;
      data_in <= ptr_deref_49_data_0 & ptr_deref_77_data_0 & ptr_deref_135_data_0 & ptr_deref_157_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 7,
        data_width => 16,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(6 downto 0),
          mdata => memory_space_1_sr_data(15 downto 0),
          mtag => memory_space_1_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 4,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : ptr_deref_302_store_0 ptr_deref_324_store_0 ptr_deref_223_store_0 ptr_deref_251_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_302_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_324_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_223_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_251_store_0_req_0;
      ptr_deref_302_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_324_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_223_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_251_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_302_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_324_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_223_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_251_store_0_req_1;
      ptr_deref_302_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_324_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_223_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_251_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      StoreGroup4_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup4_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup4_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup4_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup4_gI: SplitGuardInterface generic map(name => "StoreGroup4_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_302_word_address_0 & ptr_deref_324_word_address_0 & ptr_deref_223_word_address_0 & ptr_deref_251_word_address_0;
      data_in <= ptr_deref_302_data_0 & ptr_deref_324_data_0 & ptr_deref_223_data_0 & ptr_deref_251_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup4 Req ", addr_width => 7,
        data_width => 16,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(6 downto 0),
          mdata => memory_space_2_sr_data(15 downto 0),
          mtag => memory_space_2_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup4 Complete ",
          num_reqs => 4,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : ptr_deref_392_store_0 ptr_deref_414_store_0 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(1 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_392_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_414_store_0_req_0;
      ptr_deref_392_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_414_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_392_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_414_store_0_req_1;
      ptr_deref_392_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_414_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup5_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup5_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup5_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup5_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup5_gI: SplitGuardInterface generic map(name => "StoreGroup5_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_392_word_address_0 & ptr_deref_414_word_address_0;
      data_in <= ptr_deref_392_data_0 & ptr_deref_414_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup5 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_8_sr_req(0),
          mack => memory_space_8_sr_ack(0),
          maddr => memory_space_8_sr_addr(0 downto 0),
          mdata => memory_space_8_sr_data(15 downto 0),
          mtag => memory_space_8_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup5 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_8_sc_req(0),
          mack => memory_space_8_sc_ack(0),
          mtag => memory_space_8_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared store operator group (6) : ptr_deref_545_store_0 ptr_deref_496_store_0 ptr_deref_575_store_0 ptr_deref_624_store_0 ptr_deref_526_store_0 ptr_deref_594_store_0 
    StoreGroup6: Block -- 
      signal addr_in: std_logic_vector(41 downto 0);
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 5 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 5 downto 0);
      signal guard_vector : std_logic_vector( 5 downto 0);
      constant inBUFs : IntegerArray(5 downto 0) := (5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(5 downto 0) := (5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(5 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false);
      constant guardBuffering: IntegerArray(5 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2);
      -- 
    begin -- 
      reqL_unguarded(5) <= ptr_deref_545_store_0_req_0;
      reqL_unguarded(4) <= ptr_deref_496_store_0_req_0;
      reqL_unguarded(3) <= ptr_deref_575_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_624_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_526_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_594_store_0_req_0;
      ptr_deref_545_store_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_496_store_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_575_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_624_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_526_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_594_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(5) <= ptr_deref_545_store_0_req_1;
      reqR_unguarded(4) <= ptr_deref_496_store_0_req_1;
      reqR_unguarded(3) <= ptr_deref_575_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_624_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_526_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_594_store_0_req_1;
      ptr_deref_545_store_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_496_store_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_575_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_624_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_526_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_594_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      StoreGroup6_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup6_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup6_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup6_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup6_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup6_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup6_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup6_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup6_accessRegulator_4: access_regulator_base generic map (name => "StoreGroup6_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      StoreGroup6_accessRegulator_5: access_regulator_base generic map (name => "StoreGroup6_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      StoreGroup6_gI: SplitGuardInterface generic map(name => "StoreGroup6_gI", nreqs => 6, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_545_word_address_0 & ptr_deref_496_word_address_0 & ptr_deref_575_word_address_0 & ptr_deref_624_word_address_0 & ptr_deref_526_word_address_0 & ptr_deref_594_word_address_0;
      data_in <= ptr_deref_545_data_0 & ptr_deref_496_data_0 & ptr_deref_575_data_0 & ptr_deref_624_data_0 & ptr_deref_526_data_0 & ptr_deref_594_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup6 Req ", addr_width => 7,
        data_width => 16,
        num_reqs => 6,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(6 downto 0),
          mdata => memory_space_3_sr_data(15 downto 0),
          mtag => memory_space_3_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup6 Complete ",
          num_reqs => 6,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 6
    -- shared store operator group (7) : ptr_deref_978_store_0 
    StoreGroup7: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_978_store_0_req_0;
      ptr_deref_978_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_978_store_0_req_1;
      ptr_deref_978_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup7_gI: SplitGuardInterface generic map(name => "StoreGroup7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_978_word_address_0;
      data_in <= ptr_deref_978_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup7 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(13 downto 0),
          mdata => memory_space_4_sr_data(63 downto 0),
          mtag => memory_space_4_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup7 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 7
    -- shared inport operator group (0) : RPIPE_ConvTranspose_input_pipe_530_inst RPIPE_ConvTranspose_input_pipe_295_inst RPIPE_ConvTranspose_input_pipe_312_inst RPIPE_ConvTranspose_input_pipe_481_inst RPIPE_ConvTranspose_input_pipe_555_inst RPIPE_ConvTranspose_input_pipe_402_inst RPIPE_ConvTranspose_input_pipe_604_inst RPIPE_ConvTranspose_input_pipe_364_inst RPIPE_ConvTranspose_input_pipe_506_inst RPIPE_ConvTranspose_input_pipe_418_inst RPIPE_ConvTranspose_input_pipe_579_inst RPIPE_ConvTranspose_input_pipe_466_inst RPIPE_ConvTranspose_input_pipe_36_inst RPIPE_ConvTranspose_input_pipe_59_inst RPIPE_ConvTranspose_input_pipe_88_inst RPIPE_ConvTranspose_input_pipe_145_inst RPIPE_ConvTranspose_input_pipe_189_inst RPIPE_ConvTranspose_input_pipe_233_inst RPIPE_ConvTranspose_input_pipe_845_inst RPIPE_ConvTranspose_input_pipe_858_inst RPIPE_ConvTranspose_input_pipe_876_inst RPIPE_ConvTranspose_input_pipe_894_inst RPIPE_ConvTranspose_input_pipe_912_inst RPIPE_ConvTranspose_input_pipe_930_inst RPIPE_ConvTranspose_input_pipe_948_inst RPIPE_ConvTranspose_input_pipe_966_inst RPIPE_ConvTranspose_input_pipe_1052_inst RPIPE_ConvTranspose_input_pipe_1065_inst RPIPE_ConvTranspose_input_pipe_1083_inst RPIPE_ConvTranspose_input_pipe_1101_inst RPIPE_ConvTranspose_input_pipe_1119_inst RPIPE_ConvTranspose_input_pipe_1137_inst RPIPE_ConvTranspose_input_pipe_1155_inst RPIPE_ConvTranspose_input_pipe_1173_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(271 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 33 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 33 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 33 downto 0);
      signal guard_vector : std_logic_vector( 33 downto 0);
      constant outBUFs : IntegerArray(33 downto 0) := (33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(33 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false);
      constant guardBuffering: IntegerArray(33 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2);
      -- 
    begin -- 
      reqL_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_530_inst_req_0;
      reqL_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_295_inst_req_0;
      reqL_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_312_inst_req_0;
      reqL_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_481_inst_req_0;
      reqL_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_555_inst_req_0;
      reqL_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_402_inst_req_0;
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_604_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_364_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_506_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_418_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_579_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_466_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_36_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_59_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_88_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_145_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_189_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_233_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_845_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_858_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_876_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_894_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_912_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_930_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_948_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_966_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_1052_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_1065_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_1083_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_1101_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_1119_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_1137_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_1155_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_1173_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_530_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_295_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_312_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_481_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_555_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_402_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_604_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_364_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_506_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_418_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_579_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_466_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_36_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_59_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_88_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_145_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_189_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_233_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_845_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_858_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_876_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_894_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_912_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_930_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_948_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_966_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_1052_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_1065_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_1083_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_1101_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_1119_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_1137_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_1155_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_1173_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_530_inst_req_1;
      reqR_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_295_inst_req_1;
      reqR_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_312_inst_req_1;
      reqR_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_481_inst_req_1;
      reqR_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_555_inst_req_1;
      reqR_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_402_inst_req_1;
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_604_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_364_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_506_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_418_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_579_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_466_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_36_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_59_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_88_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_145_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_189_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_233_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_845_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_858_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_876_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_894_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_912_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_930_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_948_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_966_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_1052_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_1065_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_1083_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_1101_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_1119_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_1137_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_1155_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_1173_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_530_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_295_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_312_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_481_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_555_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_402_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_604_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_364_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_506_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_418_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_579_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_466_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_36_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_59_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_88_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_145_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_189_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_233_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_845_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_858_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_876_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_894_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_912_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_930_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_948_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_966_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_1052_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_1065_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_1083_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_1101_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_1119_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_1137_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_1155_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_1173_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      call110_531 <= data_out(271 downto 264);
      call43_296 <= data_out(263 downto 256);
      call54_313 <= data_out(255 downto 248);
      call101_482 <= data_out(247 downto 240);
      call115_556 <= data_out(239 downto 232);
      call81_403 <= data_out(231 downto 224);
      call124_605 <= data_out(223 downto 216);
      call70303_365 <= data_out(215 downto 208);
      call106_507 <= data_out(207 downto 200);
      call70_419 <= data_out(199 downto 192);
      call119_580 <= data_out(191 downto 184);
      call97_467 <= data_out(183 downto 176);
      call_37 <= data_out(175 downto 168);
      call2_60 <= data_out(167 downto 160);
      call10317_89 <= data_out(159 downto 152);
      call19_146 <= data_out(151 downto 144);
      call10_190 <= data_out(143 downto 136);
      call32_234 <= data_out(135 downto 128);
      call155_846 <= data_out(127 downto 120);
      call159_859 <= data_out(119 downto 112);
      call165_877 <= data_out(111 downto 104);
      call171_895 <= data_out(103 downto 96);
      call177_913 <= data_out(95 downto 88);
      call183_931 <= data_out(87 downto 80);
      call189_949 <= data_out(79 downto 72);
      call195_967 <= data_out(71 downto 64);
      call216_1053 <= data_out(63 downto 56);
      call220_1066 <= data_out(55 downto 48);
      call226_1084 <= data_out(47 downto 40);
      call232_1102 <= data_out(39 downto 32);
      call238_1120 <= data_out(31 downto 24);
      call244_1138 <= data_out(23 downto 16);
      call250_1156 <= data_out(15 downto 8);
      call256_1174 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_0_gI", nreqs => 34, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_0", data_width => 8,  num_reqs => 34,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end testConfigure_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(31 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(31 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_4124_start: Boolean;
  signal timer_CP_4124_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_1367_load_0_req_0 : boolean;
  signal LOAD_count_1367_load_0_ack_0 : boolean;
  signal LOAD_count_1367_load_0_req_1 : boolean;
  signal LOAD_count_1367_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_4124_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= c_buffer;
  c <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_4124_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_4124_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_4124_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_4124: Block -- control-path 
    signal timer_CP_4124_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_4124_elements(0) <= timer_CP_4124_start;
    timer_CP_4124_symbol <= timer_CP_4124_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_1368/$entry
      -- CP-element group 0: 	 assign_stmt_1368/LOAD_count_1367_sample_start_
      -- CP-element group 0: 	 assign_stmt_1368/LOAD_count_1367_update_start_
      -- CP-element group 0: 	 assign_stmt_1368/LOAD_count_1367_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_1368/LOAD_count_1367_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_1368/LOAD_count_1367_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1368/LOAD_count_1367_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_1368/LOAD_count_1367_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_1368/LOAD_count_1367_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_1368/LOAD_count_1367_Update/$entry
      -- CP-element group 0: 	 assign_stmt_1368/LOAD_count_1367_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_1368/LOAD_count_1367_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_1368/LOAD_count_1367_Update/word_access_complete/word_0/cr
      -- 
    rr_4145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_4124_elements(0), ack => LOAD_count_1367_load_0_req_0); -- 
    cr_4156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_4124_elements(0), ack => LOAD_count_1367_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_1368/LOAD_count_1367_sample_completed_
      -- CP-element group 1: 	 assign_stmt_1368/LOAD_count_1367_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1368/LOAD_count_1367_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_1368/LOAD_count_1367_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_1368/LOAD_count_1367_Sample/word_access_start/word_0/ra
      -- 
    ra_4146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_1367_load_0_ack_0, ack => timer_CP_4124_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_1368/$exit
      -- CP-element group 2: 	 assign_stmt_1368/LOAD_count_1367_update_completed_
      -- CP-element group 2: 	 assign_stmt_1368/LOAD_count_1367_Update/$exit
      -- CP-element group 2: 	 assign_stmt_1368/LOAD_count_1367_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_1368/LOAD_count_1367_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_1368/LOAD_count_1367_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_1368/LOAD_count_1367_Update/LOAD_count_1367_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_1368/LOAD_count_1367_Update/LOAD_count_1367_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_1368/LOAD_count_1367_Update/LOAD_count_1367_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_1368/LOAD_count_1367_Update/LOAD_count_1367_Merge/merge_ack
      -- 
    ca_4157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_1367_load_0_ack_1, ack => timer_CP_4124_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_1367_data_0 : std_logic_vector(31 downto 0);
    signal LOAD_count_1367_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_1367_word_address_0 <= "0";
    -- equivalence LOAD_count_1367_gather_scatter
    process(LOAD_count_1367_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_1367_data_0;
      ov(31 downto 0) := iv;
      c_buffer <= ov(31 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_1367_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_1367_load_0_req_0;
      LOAD_count_1367_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_1367_load_0_req_1;
      LOAD_count_1367_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_1367_word_address_0;
      LOAD_count_1367_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(4 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(4 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(34 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(104 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(4 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(79 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(14 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(4 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(4 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(34 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(104 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(4 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(79 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(14 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(5 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(5 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(41 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(125 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(5 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(5 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(95 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(17 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_4_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_4_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_4_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_4_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_4_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_4_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_4_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_5
  signal memory_space_5_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_5_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_5_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_5_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_5_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_5_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_5_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_5_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_6
  signal memory_space_6_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_6_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_6_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_6_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_6_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_6_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_6_sr_addr : std_logic_vector(69 downto 0);
  signal memory_space_6_sr_data : std_logic_vector(319 downto 0);
  signal memory_space_6_sr_tag : std_logic_vector(94 downto 0);
  signal memory_space_6_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_6_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_6_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_7
  signal memory_space_7_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_7_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_7_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_7_lr_tag : std_logic_vector(79 downto 0);
  signal memory_space_7_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_7_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_7_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_7_lc_tag :  std_logic_vector(7 downto 0);
  signal memory_space_7_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_7_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_7_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_8
  signal memory_space_8_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_8_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_8_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_8_lr_tag : std_logic_vector(79 downto 0);
  signal memory_space_8_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_8_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_8_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_8_lc_tag :  std_logic_vector(7 downto 0);
  signal memory_space_8_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_8_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_8_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_sc_tag :  std_logic_vector(1 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_call_acks : in   std_logic_vector(0 downto 0);
      testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
      testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_return_acks : in   std_logic_vector(0 downto 0);
      testConfigure_return_data : in   std_logic_vector(15 downto 0);
      testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(31 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_call_acks : in   std_logic_vector(0 downto 0);
      sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
      sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_return_acks : in   std_logic_vector(0 downto 0);
      sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module sendOutput
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendOutput
  signal sendOutput_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendOutput_tag_out   : std_logic_vector(1 downto 0);
  signal sendOutput_start_req : std_logic;
  signal sendOutput_start_ack : std_logic;
  signal sendOutput_fin_req   : std_logic;
  signal sendOutput_fin_ack : std_logic;
  -- caller side aggregated signals for module sendOutput
  signal sendOutput_call_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_call_acks: std_logic_vector(0 downto 0);
  signal sendOutput_return_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_return_acks: std_logic_vector(0 downto 0);
  signal sendOutput_call_tag: std_logic_vector(0 downto 0);
  signal sendOutput_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module testConfigure
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module testConfigure
  signal testConfigure_ret_val_x_x :  std_logic_vector(15 downto 0);
  signal testConfigure_out_args   : std_logic_vector(15 downto 0);
  signal testConfigure_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal testConfigure_tag_out   : std_logic_vector(1 downto 0);
  signal testConfigure_start_req : std_logic;
  signal testConfigure_start_ack : std_logic;
  signal testConfigure_fin_req   : std_logic;
  signal testConfigure_fin_ack : std_logic;
  -- caller side aggregated signals for module testConfigure
  signal testConfigure_call_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_call_acks: std_logic_vector(0 downto 0);
  signal testConfigure_return_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_return_acks: std_logic_vector(0 downto 0);
  signal testConfigure_call_tag: std_logic_vector(0 downto 0);
  signal testConfigure_return_data: std_logic_vector(15 downto 0);
  signal testConfigure_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(31 downto 0);
  signal timer_out_args   : std_logic_vector(31 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(31 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_start
  signal Block2_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_start
  signal Block3_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(15 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(15 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(15 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(15 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(15 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(15 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      testConfigure_call_reqs => testConfigure_call_reqs(0 downto 0),
      testConfigure_call_acks => testConfigure_call_acks(0 downto 0),
      testConfigure_call_tag => testConfigure_call_tag(0 downto 0),
      testConfigure_return_reqs => testConfigure_return_reqs(0 downto 0),
      testConfigure_return_acks => testConfigure_return_acks(0 downto 0),
      testConfigure_return_data => testConfigure_return_data(15 downto 0),
      testConfigure_return_tag => testConfigure_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(31 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      sendOutput_call_reqs => sendOutput_call_reqs(0 downto 0),
      sendOutput_call_acks => sendOutput_call_acks(0 downto 0),
      sendOutput_call_tag => sendOutput_call_tag(0 downto 0),
      sendOutput_return_reqs => sendOutput_return_reqs(0 downto 0),
      sendOutput_return_acks => sendOutput_return_acks(0 downto 0),
      sendOutput_return_tag => sendOutput_return_tag(0 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(3 downto 3),
      memory_space_1_lr_ack => memory_space_1_lr_ack(3 downto 3),
      memory_space_1_lr_addr => memory_space_1_lr_addr(27 downto 21),
      memory_space_1_lr_tag => memory_space_1_lr_tag(83 downto 63),
      memory_space_1_lc_req => memory_space_1_lc_req(3 downto 3),
      memory_space_1_lc_ack => memory_space_1_lc_ack(3 downto 3),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 48),
      memory_space_1_lc_tag => memory_space_1_lc_tag(11 downto 9),
      memory_space_2_lr_req => memory_space_2_lr_req(3 downto 3),
      memory_space_2_lr_ack => memory_space_2_lr_ack(3 downto 3),
      memory_space_2_lr_addr => memory_space_2_lr_addr(27 downto 21),
      memory_space_2_lr_tag => memory_space_2_lr_tag(83 downto 63),
      memory_space_2_lc_req => memory_space_2_lc_req(3 downto 3),
      memory_space_2_lc_ack => memory_space_2_lc_ack(3 downto 3),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 48),
      memory_space_2_lc_tag => memory_space_2_lc_tag(11 downto 9),
      memory_space_3_lr_req => memory_space_3_lr_req(3 downto 3),
      memory_space_3_lr_ack => memory_space_3_lr_ack(3 downto 3),
      memory_space_3_lr_addr => memory_space_3_lr_addr(27 downto 21),
      memory_space_3_lr_tag => memory_space_3_lr_tag(83 downto 63),
      memory_space_3_lc_req => memory_space_3_lc_req(3 downto 3),
      memory_space_3_lc_ack => memory_space_3_lc_ack(3 downto 3),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 48),
      memory_space_3_lc_tag => memory_space_3_lc_tag(11 downto 9),
      memory_space_4_lr_req => memory_space_4_lr_req(3 downto 3),
      memory_space_4_lr_ack => memory_space_4_lr_ack(3 downto 3),
      memory_space_4_lr_addr => memory_space_4_lr_addr(55 downto 42),
      memory_space_4_lr_tag => memory_space_4_lr_tag(75 downto 57),
      memory_space_4_lc_req => memory_space_4_lc_req(3 downto 3),
      memory_space_4_lc_ack => memory_space_4_lc_ack(3 downto 3),
      memory_space_4_lc_data => memory_space_4_lc_data(255 downto 192),
      memory_space_4_lc_tag => memory_space_4_lc_tag(3 downto 3),
      memory_space_7_lr_req => memory_space_7_lr_req(3 downto 3),
      memory_space_7_lr_ack => memory_space_7_lr_ack(3 downto 3),
      memory_space_7_lr_addr => memory_space_7_lr_addr(3 downto 3),
      memory_space_7_lr_tag => memory_space_7_lr_tag(79 downto 60),
      memory_space_7_lc_req => memory_space_7_lc_req(3 downto 3),
      memory_space_7_lc_ack => memory_space_7_lc_ack(3 downto 3),
      memory_space_7_lc_data => memory_space_7_lc_data(63 downto 48),
      memory_space_7_lc_tag => memory_space_7_lc_tag(7 downto 6),
      memory_space_8_lr_req => memory_space_8_lr_req(3 downto 3),
      memory_space_8_lr_ack => memory_space_8_lr_ack(3 downto 3),
      memory_space_8_lr_addr => memory_space_8_lr_addr(3 downto 3),
      memory_space_8_lr_tag => memory_space_8_lr_tag(79 downto 60),
      memory_space_8_lc_req => memory_space_8_lc_req(3 downto 3),
      memory_space_8_lc_ack => memory_space_8_lc_ack(3 downto 3),
      memory_space_8_lc_data => memory_space_8_lc_data(63 downto 48),
      memory_space_8_lc_tag => memory_space_8_lc_tag(7 downto 6),
      memory_space_6_sr_req => memory_space_6_sr_req(3 downto 3),
      memory_space_6_sr_ack => memory_space_6_sr_ack(3 downto 3),
      memory_space_6_sr_addr => memory_space_6_sr_addr(55 downto 42),
      memory_space_6_sr_data => memory_space_6_sr_data(255 downto 192),
      memory_space_6_sr_tag => memory_space_6_sr_tag(75 downto 57),
      memory_space_6_sc_req => memory_space_6_sc_req(3 downto 3),
      memory_space_6_sc_ack => memory_space_6_sc_ack(3 downto 3),
      memory_space_6_sc_tag => memory_space_6_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(20 downto 14),
      memory_space_1_lr_tag => memory_space_1_lr_tag(62 downto 42),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(47 downto 32),
      memory_space_1_lc_tag => memory_space_1_lc_tag(8 downto 6),
      memory_space_2_lr_req => memory_space_2_lr_req(2 downto 2),
      memory_space_2_lr_ack => memory_space_2_lr_ack(2 downto 2),
      memory_space_2_lr_addr => memory_space_2_lr_addr(20 downto 14),
      memory_space_2_lr_tag => memory_space_2_lr_tag(62 downto 42),
      memory_space_2_lc_req => memory_space_2_lc_req(2 downto 2),
      memory_space_2_lc_ack => memory_space_2_lc_ack(2 downto 2),
      memory_space_2_lc_data => memory_space_2_lc_data(47 downto 32),
      memory_space_2_lc_tag => memory_space_2_lc_tag(8 downto 6),
      memory_space_3_lr_req => memory_space_3_lr_req(2 downto 2),
      memory_space_3_lr_ack => memory_space_3_lr_ack(2 downto 2),
      memory_space_3_lr_addr => memory_space_3_lr_addr(20 downto 14),
      memory_space_3_lr_tag => memory_space_3_lr_tag(62 downto 42),
      memory_space_3_lc_req => memory_space_3_lc_req(2 downto 2),
      memory_space_3_lc_ack => memory_space_3_lc_ack(2 downto 2),
      memory_space_3_lc_data => memory_space_3_lc_data(47 downto 32),
      memory_space_3_lc_tag => memory_space_3_lc_tag(8 downto 6),
      memory_space_4_lr_req => memory_space_4_lr_req(2 downto 2),
      memory_space_4_lr_ack => memory_space_4_lr_ack(2 downto 2),
      memory_space_4_lr_addr => memory_space_4_lr_addr(41 downto 28),
      memory_space_4_lr_tag => memory_space_4_lr_tag(56 downto 38),
      memory_space_4_lc_req => memory_space_4_lc_req(2 downto 2),
      memory_space_4_lc_ack => memory_space_4_lc_ack(2 downto 2),
      memory_space_4_lc_data => memory_space_4_lc_data(191 downto 128),
      memory_space_4_lc_tag => memory_space_4_lc_tag(2 downto 2),
      memory_space_7_lr_req => memory_space_7_lr_req(2 downto 2),
      memory_space_7_lr_ack => memory_space_7_lr_ack(2 downto 2),
      memory_space_7_lr_addr => memory_space_7_lr_addr(2 downto 2),
      memory_space_7_lr_tag => memory_space_7_lr_tag(59 downto 40),
      memory_space_7_lc_req => memory_space_7_lc_req(2 downto 2),
      memory_space_7_lc_ack => memory_space_7_lc_ack(2 downto 2),
      memory_space_7_lc_data => memory_space_7_lc_data(47 downto 32),
      memory_space_7_lc_tag => memory_space_7_lc_tag(5 downto 4),
      memory_space_8_lr_req => memory_space_8_lr_req(2 downto 2),
      memory_space_8_lr_ack => memory_space_8_lr_ack(2 downto 2),
      memory_space_8_lr_addr => memory_space_8_lr_addr(2 downto 2),
      memory_space_8_lr_tag => memory_space_8_lr_tag(59 downto 40),
      memory_space_8_lc_req => memory_space_8_lc_req(2 downto 2),
      memory_space_8_lc_ack => memory_space_8_lc_ack(2 downto 2),
      memory_space_8_lc_data => memory_space_8_lc_data(47 downto 32),
      memory_space_8_lc_tag => memory_space_8_lc_tag(5 downto 4),
      memory_space_6_sr_req => memory_space_6_sr_req(2 downto 2),
      memory_space_6_sr_ack => memory_space_6_sr_ack(2 downto 2),
      memory_space_6_sr_addr => memory_space_6_sr_addr(41 downto 28),
      memory_space_6_sr_data => memory_space_6_sr_data(191 downto 128),
      memory_space_6_sr_tag => memory_space_6_sr_tag(56 downto 38),
      memory_space_6_sc_req => memory_space_6_sc_req(2 downto 2),
      memory_space_6_sc_ack => memory_space_6_sc_ack(2 downto 2),
      memory_space_6_sc_tag => memory_space_6_sc_tag(2 downto 2),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(15 downto 0),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 7),
      memory_space_1_lr_tag => memory_space_1_lr_tag(41 downto 21),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(31 downto 16),
      memory_space_1_lc_tag => memory_space_1_lc_tag(5 downto 3),
      memory_space_2_lr_req => memory_space_2_lr_req(1 downto 1),
      memory_space_2_lr_ack => memory_space_2_lr_ack(1 downto 1),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 7),
      memory_space_2_lr_tag => memory_space_2_lr_tag(41 downto 21),
      memory_space_2_lc_req => memory_space_2_lc_req(1 downto 1),
      memory_space_2_lc_ack => memory_space_2_lc_ack(1 downto 1),
      memory_space_2_lc_data => memory_space_2_lc_data(31 downto 16),
      memory_space_2_lc_tag => memory_space_2_lc_tag(5 downto 3),
      memory_space_3_lr_req => memory_space_3_lr_req(1 downto 1),
      memory_space_3_lr_ack => memory_space_3_lr_ack(1 downto 1),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 7),
      memory_space_3_lr_tag => memory_space_3_lr_tag(41 downto 21),
      memory_space_3_lc_req => memory_space_3_lc_req(1 downto 1),
      memory_space_3_lc_ack => memory_space_3_lc_ack(1 downto 1),
      memory_space_3_lc_data => memory_space_3_lc_data(31 downto 16),
      memory_space_3_lc_tag => memory_space_3_lc_tag(5 downto 3),
      memory_space_4_lr_req => memory_space_4_lr_req(1 downto 1),
      memory_space_4_lr_ack => memory_space_4_lr_ack(1 downto 1),
      memory_space_4_lr_addr => memory_space_4_lr_addr(27 downto 14),
      memory_space_4_lr_tag => memory_space_4_lr_tag(37 downto 19),
      memory_space_4_lc_req => memory_space_4_lc_req(1 downto 1),
      memory_space_4_lc_ack => memory_space_4_lc_ack(1 downto 1),
      memory_space_4_lc_data => memory_space_4_lc_data(127 downto 64),
      memory_space_4_lc_tag => memory_space_4_lc_tag(1 downto 1),
      memory_space_7_lr_req => memory_space_7_lr_req(1 downto 1),
      memory_space_7_lr_ack => memory_space_7_lr_ack(1 downto 1),
      memory_space_7_lr_addr => memory_space_7_lr_addr(1 downto 1),
      memory_space_7_lr_tag => memory_space_7_lr_tag(39 downto 20),
      memory_space_7_lc_req => memory_space_7_lc_req(1 downto 1),
      memory_space_7_lc_ack => memory_space_7_lc_ack(1 downto 1),
      memory_space_7_lc_data => memory_space_7_lc_data(31 downto 16),
      memory_space_7_lc_tag => memory_space_7_lc_tag(3 downto 2),
      memory_space_8_lr_req => memory_space_8_lr_req(1 downto 1),
      memory_space_8_lr_ack => memory_space_8_lr_ack(1 downto 1),
      memory_space_8_lr_addr => memory_space_8_lr_addr(1 downto 1),
      memory_space_8_lr_tag => memory_space_8_lr_tag(39 downto 20),
      memory_space_8_lc_req => memory_space_8_lc_req(1 downto 1),
      memory_space_8_lc_ack => memory_space_8_lc_ack(1 downto 1),
      memory_space_8_lc_data => memory_space_8_lc_data(31 downto 16),
      memory_space_8_lc_tag => memory_space_8_lc_tag(3 downto 2),
      memory_space_6_sr_req => memory_space_6_sr_req(1 downto 1),
      memory_space_6_sr_ack => memory_space_6_sr_ack(1 downto 1),
      memory_space_6_sr_addr => memory_space_6_sr_addr(27 downto 14),
      memory_space_6_sr_data => memory_space_6_sr_data(127 downto 64),
      memory_space_6_sr_tag => memory_space_6_sr_tag(37 downto 19),
      memory_space_6_sc_req => memory_space_6_sc_req(1 downto 1),
      memory_space_6_sc_ack => memory_space_6_sc_ack(1 downto 1),
      memory_space_6_sc_tag => memory_space_6_sc_tag(1 downto 1),
      Block2_start_pipe_read_req => Block2_start_pipe_read_req(0 downto 0),
      Block2_start_pipe_read_ack => Block2_start_pipe_read_ack(0 downto 0),
      Block2_start_pipe_read_data => Block2_start_pipe_read_data(15 downto 0),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(6 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(20 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(15 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(6 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(20 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(15 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(2 downto 0),
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(6 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(20 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(15 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(2 downto 0),
      memory_space_4_lr_req => memory_space_4_lr_req(0 downto 0),
      memory_space_4_lr_ack => memory_space_4_lr_ack(0 downto 0),
      memory_space_4_lr_addr => memory_space_4_lr_addr(13 downto 0),
      memory_space_4_lr_tag => memory_space_4_lr_tag(18 downto 0),
      memory_space_4_lc_req => memory_space_4_lc_req(0 downto 0),
      memory_space_4_lc_ack => memory_space_4_lc_ack(0 downto 0),
      memory_space_4_lc_data => memory_space_4_lc_data(63 downto 0),
      memory_space_4_lc_tag => memory_space_4_lc_tag(0 downto 0),
      memory_space_7_lr_req => memory_space_7_lr_req(0 downto 0),
      memory_space_7_lr_ack => memory_space_7_lr_ack(0 downto 0),
      memory_space_7_lr_addr => memory_space_7_lr_addr(0 downto 0),
      memory_space_7_lr_tag => memory_space_7_lr_tag(19 downto 0),
      memory_space_7_lc_req => memory_space_7_lc_req(0 downto 0),
      memory_space_7_lc_ack => memory_space_7_lc_ack(0 downto 0),
      memory_space_7_lc_data => memory_space_7_lc_data(15 downto 0),
      memory_space_7_lc_tag => memory_space_7_lc_tag(1 downto 0),
      memory_space_8_lr_req => memory_space_8_lr_req(0 downto 0),
      memory_space_8_lr_ack => memory_space_8_lr_ack(0 downto 0),
      memory_space_8_lr_addr => memory_space_8_lr_addr(0 downto 0),
      memory_space_8_lr_tag => memory_space_8_lr_tag(19 downto 0),
      memory_space_8_lc_req => memory_space_8_lc_req(0 downto 0),
      memory_space_8_lc_ack => memory_space_8_lc_ack(0 downto 0),
      memory_space_8_lc_data => memory_space_8_lc_data(15 downto 0),
      memory_space_8_lc_tag => memory_space_8_lc_tag(1 downto 0),
      memory_space_6_sr_req => memory_space_6_sr_req(0 downto 0),
      memory_space_6_sr_ack => memory_space_6_sr_ack(0 downto 0),
      memory_space_6_sr_addr => memory_space_6_sr_addr(13 downto 0),
      memory_space_6_sr_data => memory_space_6_sr_data(63 downto 0),
      memory_space_6_sr_tag => memory_space_6_sr_tag(18 downto 0),
      memory_space_6_sc_req => memory_space_6_sc_req(0 downto 0),
      memory_space_6_sc_ack => memory_space_6_sc_ack(0 downto 0),
      memory_space_6_sc_tag => memory_space_6_sc_tag(0 downto 0),
      Block3_start_pipe_read_req => Block3_start_pipe_read_req(0 downto 0),
      Block3_start_pipe_read_ack => Block3_start_pipe_read_ack(0 downto 0),
      Block3_start_pipe_read_data => Block3_start_pipe_read_data(15 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module sendOutput
  -- call arbiter for module sendOutput
  sendOutput_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendOutput_call_reqs,
      call_acks => sendOutput_call_acks,
      return_reqs => sendOutput_return_reqs,
      return_acks => sendOutput_return_acks,
      call_tag  => sendOutput_call_tag,
      return_tag  => sendOutput_return_tag,
      call_mtag => sendOutput_tag_in,
      return_mtag => sendOutput_tag_out,
      call_mreq => sendOutput_start_req,
      call_mack => sendOutput_start_ack,
      return_mreq => sendOutput_fin_req,
      return_mack => sendOutput_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  sendOutput_instance:sendOutput-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendOutput_start_req,
      start_ack => sendOutput_start_ack,
      fin_req => sendOutput_fin_req,
      fin_ack => sendOutput_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(4 downto 4),
      memory_space_3_lr_ack => memory_space_3_lr_ack(4 downto 4),
      memory_space_3_lr_addr => memory_space_3_lr_addr(34 downto 28),
      memory_space_3_lr_tag => memory_space_3_lr_tag(104 downto 84),
      memory_space_3_lc_req => memory_space_3_lc_req(4 downto 4),
      memory_space_3_lc_ack => memory_space_3_lc_ack(4 downto 4),
      memory_space_3_lc_data => memory_space_3_lc_data(79 downto 64),
      memory_space_3_lc_tag => memory_space_3_lc_tag(14 downto 12),
      memory_space_6_lr_req => memory_space_6_lr_req(0 downto 0),
      memory_space_6_lr_ack => memory_space_6_lr_ack(0 downto 0),
      memory_space_6_lr_addr => memory_space_6_lr_addr(13 downto 0),
      memory_space_6_lr_tag => memory_space_6_lr_tag(18 downto 0),
      memory_space_6_lc_req => memory_space_6_lc_req(0 downto 0),
      memory_space_6_lc_ack => memory_space_6_lc_ack(0 downto 0),
      memory_space_6_lc_data => memory_space_6_lc_data(63 downto 0),
      memory_space_6_lc_tag => memory_space_6_lc_tag(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      tag_in => sendOutput_tag_in,
      tag_out => sendOutput_tag_out-- 
    ); -- 
  -- module testConfigure
  testConfigure_out_args <= testConfigure_ret_val_x_x ;
  -- call arbiter for module testConfigure
  testConfigure_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 16,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => testConfigure_call_reqs,
      call_acks => testConfigure_call_acks,
      return_reqs => testConfigure_return_reqs,
      return_acks => testConfigure_return_acks,
      call_tag  => testConfigure_call_tag,
      return_tag  => testConfigure_return_tag,
      call_mtag => testConfigure_tag_in,
      return_mtag => testConfigure_tag_out,
      return_data =>testConfigure_return_data,
      call_mreq => testConfigure_start_req,
      call_mack => testConfigure_start_ack,
      return_mreq => testConfigure_fin_req,
      return_mack => testConfigure_fin_ack,
      return_mdata => testConfigure_out_args,
      clk => clk, 
      reset => reset --
    ); --
  testConfigure_instance:testConfigure-- 
    generic map(tag_length => 2)
    port map(-- 
      ret_val_x_x => testConfigure_ret_val_x_x,
      start_req => testConfigure_start_req,
      start_ack => testConfigure_start_ack,
      fin_req => testConfigure_fin_req,
      fin_ack => testConfigure_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(4 downto 4),
      memory_space_1_lr_ack => memory_space_1_lr_ack(4 downto 4),
      memory_space_1_lr_addr => memory_space_1_lr_addr(34 downto 28),
      memory_space_1_lr_tag => memory_space_1_lr_tag(104 downto 84),
      memory_space_1_lc_req => memory_space_1_lc_req(4 downto 4),
      memory_space_1_lc_ack => memory_space_1_lc_ack(4 downto 4),
      memory_space_1_lc_data => memory_space_1_lc_data(79 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(14 downto 12),
      memory_space_2_lr_req => memory_space_2_lr_req(4 downto 4),
      memory_space_2_lr_ack => memory_space_2_lr_ack(4 downto 4),
      memory_space_2_lr_addr => memory_space_2_lr_addr(34 downto 28),
      memory_space_2_lr_tag => memory_space_2_lr_tag(104 downto 84),
      memory_space_2_lc_req => memory_space_2_lc_req(4 downto 4),
      memory_space_2_lc_ack => memory_space_2_lc_ack(4 downto 4),
      memory_space_2_lc_data => memory_space_2_lc_data(79 downto 64),
      memory_space_2_lc_tag => memory_space_2_lc_tag(14 downto 12),
      memory_space_3_lr_req => memory_space_3_lr_req(5 downto 5),
      memory_space_3_lr_ack => memory_space_3_lr_ack(5 downto 5),
      memory_space_3_lr_addr => memory_space_3_lr_addr(41 downto 35),
      memory_space_3_lr_tag => memory_space_3_lr_tag(125 downto 105),
      memory_space_3_lc_req => memory_space_3_lc_req(5 downto 5),
      memory_space_3_lc_ack => memory_space_3_lc_ack(5 downto 5),
      memory_space_3_lc_data => memory_space_3_lc_data(95 downto 80),
      memory_space_3_lc_tag => memory_space_3_lc_tag(17 downto 15),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(6 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(15 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(20 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(2 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(6 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(15 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(20 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(2 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(6 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(15 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(20 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(2 downto 0),
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(13 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(63 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(18 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(0 downto 0),
      memory_space_5_sr_req => memory_space_5_sr_req(0 downto 0),
      memory_space_5_sr_ack => memory_space_5_sr_ack(0 downto 0),
      memory_space_5_sr_addr => memory_space_5_sr_addr(10 downto 0),
      memory_space_5_sr_data => memory_space_5_sr_data(63 downto 0),
      memory_space_5_sr_tag => memory_space_5_sr_tag(0 downto 0),
      memory_space_5_sc_req => memory_space_5_sc_req(0 downto 0),
      memory_space_5_sc_ack => memory_space_5_sc_ack(0 downto 0),
      memory_space_5_sc_tag => memory_space_5_sc_tag(0 downto 0),
      memory_space_6_sr_req => memory_space_6_sr_req(4 downto 4),
      memory_space_6_sr_ack => memory_space_6_sr_ack(4 downto 4),
      memory_space_6_sr_addr => memory_space_6_sr_addr(69 downto 56),
      memory_space_6_sr_data => memory_space_6_sr_data(319 downto 256),
      memory_space_6_sr_tag => memory_space_6_sr_tag(94 downto 76),
      memory_space_6_sc_req => memory_space_6_sc_req(4 downto 4),
      memory_space_6_sc_ack => memory_space_6_sc_ack(4 downto 4),
      memory_space_6_sc_tag => memory_space_6_sc_tag(4 downto 4),
      memory_space_7_sr_req => memory_space_7_sr_req(0 downto 0),
      memory_space_7_sr_ack => memory_space_7_sr_ack(0 downto 0),
      memory_space_7_sr_addr => memory_space_7_sr_addr(0 downto 0),
      memory_space_7_sr_data => memory_space_7_sr_data(15 downto 0),
      memory_space_7_sr_tag => memory_space_7_sr_tag(19 downto 0),
      memory_space_7_sc_req => memory_space_7_sc_req(0 downto 0),
      memory_space_7_sc_ack => memory_space_7_sc_ack(0 downto 0),
      memory_space_7_sc_tag => memory_space_7_sc_tag(1 downto 0),
      memory_space_8_sr_req => memory_space_8_sr_req(0 downto 0),
      memory_space_8_sr_ack => memory_space_8_sr_ack(0 downto 0),
      memory_space_8_sr_addr => memory_space_8_sr_addr(0 downto 0),
      memory_space_8_sr_data => memory_space_8_sr_data(15 downto 0),
      memory_space_8_sr_tag => memory_space_8_sr_tag(19 downto 0),
      memory_space_8_sc_req => memory_space_8_sc_req(0 downto 0),
      memory_space_8_sc_ack => memory_space_8_sc_ack(0 downto 0),
      memory_space_8_sc_tag => memory_space_8_sc_tag(1 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      tag_in => testConfigure_tag_in,
      tag_out => testConfigure_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(0 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(0 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(31 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  dummyROM_memory_space_0: dummy_read_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 5,
      num_stores => 1,
      addr_width => 7,
      data_width => 16,
      tag_width => 3,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 5,
      num_stores => 1,
      addr_width => 7,
      data_width => 16,
      tag_width => 3,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 6,
      num_stores => 1,
      addr_width => 7,
      data_width => 16,
      tag_width => 3,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_4: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_4",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_4_lr_addr,
      lr_req_in => memory_space_4_lr_req,
      lr_ack_out => memory_space_4_lr_ack,
      lr_tag_in => memory_space_4_lr_tag,
      lc_req_in => memory_space_4_lc_req,
      lc_ack_out => memory_space_4_lc_ack,
      lc_data_out => memory_space_4_lc_data,
      lc_tag_out => memory_space_4_lc_tag,
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_5: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_5",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_5_sr_addr,
      sr_data_in => memory_space_5_sr_data,
      sr_req_in => memory_space_5_sr_req,
      sr_ack_out => memory_space_5_sr_ack,
      sr_tag_in => memory_space_5_sr_tag,
      sc_req_in=> memory_space_5_sc_req,
      sc_ack_out => memory_space_5_sc_ack,
      sc_tag_out => memory_space_5_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_6: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_6",
      num_loads => 1,
      num_stores => 5,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_6_lr_addr,
      lr_req_in => memory_space_6_lr_req,
      lr_ack_out => memory_space_6_lr_ack,
      lr_tag_in => memory_space_6_lr_tag,
      lc_req_in => memory_space_6_lc_req,
      lc_ack_out => memory_space_6_lc_ack,
      lc_data_out => memory_space_6_lc_data,
      lc_tag_out => memory_space_6_lc_tag,
      sr_addr_in => memory_space_6_sr_addr,
      sr_data_in => memory_space_6_sr_data,
      sr_req_in => memory_space_6_sr_req,
      sr_ack_out => memory_space_6_sr_ack,
      sr_tag_in => memory_space_6_sr_tag,
      sc_req_in=> memory_space_6_sc_req,
      sc_ack_out => memory_space_6_sc_ack,
      sc_tag_out => memory_space_6_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_7: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_7",
      num_loads => 4,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_7_lr_addr,
      lr_req_in => memory_space_7_lr_req,
      lr_ack_out => memory_space_7_lr_ack,
      lr_tag_in => memory_space_7_lr_tag,
      lc_req_in => memory_space_7_lc_req,
      lc_ack_out => memory_space_7_lc_ack,
      lc_data_out => memory_space_7_lc_data,
      lc_tag_out => memory_space_7_lc_tag,
      sr_addr_in => memory_space_7_sr_addr,
      sr_data_in => memory_space_7_sr_data,
      sr_req_in => memory_space_7_sr_req,
      sr_ack_out => memory_space_7_sr_ack,
      sr_tag_in => memory_space_7_sr_tag,
      sc_req_in=> memory_space_7_sc_req,
      sc_ack_out => memory_space_7_sc_ack,
      sc_tag_out => memory_space_7_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_8: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_8",
      num_loads => 4,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_8_lr_addr,
      lr_req_in => memory_space_8_lr_req,
      lr_ack_out => memory_space_8_lr_ack,
      lr_tag_in => memory_space_8_lr_tag,
      lc_req_in => memory_space_8_lc_req,
      lc_ack_out => memory_space_8_lc_ack,
      lc_data_out => memory_space_8_lc_data,
      lc_tag_out => memory_space_8_lc_tag,
      sr_addr_in => memory_space_8_sr_addr,
      sr_data_in => memory_space_8_sr_data,
      sr_req_in => memory_space_8_sr_req,
      sr_ack_out => memory_space_8_sr_ack,
      sr_tag_in => memory_space_8_sr_tag,
      sc_req_in=> memory_space_8_sc_req,
      sc_ack_out => memory_space_8_sc_ack,
      sc_tag_out => memory_space_8_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
