-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(1 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    fill_kernel_call_reqs : out  std_logic_vector(0 downto 0);
    fill_kernel_call_acks : in   std_logic_vector(0 downto 0);
    fill_kernel_call_data : out  std_logic_vector(63 downto 0);
    fill_kernel_call_tag  :  out  std_logic_vector(0 downto 0);
    fill_kernel_return_reqs : out  std_logic_vector(0 downto 0);
    fill_kernel_return_acks : in   std_logic_vector(0 downto 0);
    fill_kernel_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_call_acks : in   std_logic_vector(0 downto 0);
    sendOutput_call_data : out  std_logic_vector(31 downto 0);
    sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
    sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_return_acks : in   std_logic_vector(0 downto 0);
    sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_814_start: Boolean;
  signal convTranspose_CP_814_symbol: Boolean;
  -- volatile/operator module components. 
  component fill_kernel is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(63 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(11 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_ConvTranspose_input_pipe_587_inst_ack_0 : boolean;
  signal ptr_deref_1219_store_0_ack_1 : boolean;
  signal type_cast_566_inst_req_1 : boolean;
  signal type_cast_291_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_273_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_287_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_574_inst_req_0 : boolean;
  signal type_cast_291_inst_ack_0 : boolean;
  signal type_cast_566_inst_ack_0 : boolean;
  signal addr_of_725_final_reg_ack_0 : boolean;
  signal type_cast_695_inst_req_1 : boolean;
  signal type_cast_541_inst_ack_0 : boolean;
  signal addr_of_1195_final_reg_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_728_inst_req_0 : boolean;
  signal type_cast_695_inst_ack_1 : boolean;
  signal type_cast_609_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_728_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_574_inst_ack_0 : boolean;
  signal type_cast_641_inst_req_0 : boolean;
  signal array_obj_ref_1215_index_offset_ack_1 : boolean;
  signal type_cast_578_inst_req_1 : boolean;
  signal type_cast_641_inst_ack_0 : boolean;
  signal type_cast_623_inst_ack_0 : boolean;
  signal type_cast_578_inst_ack_1 : boolean;
  signal type_cast_627_inst_req_0 : boolean;
  signal addr_of_725_final_reg_req_1 : boolean;
  signal addr_of_725_final_reg_ack_1 : boolean;
  signal type_cast_645_inst_ack_1 : boolean;
  signal type_cast_578_inst_req_0 : boolean;
  signal type_cast_605_inst_ack_1 : boolean;
  signal type_cast_605_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_299_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_728_inst_ack_1 : boolean;
  signal type_cast_303_inst_req_0 : boolean;
  signal type_cast_303_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_587_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_728_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_537_inst_req_1 : boolean;
  signal type_cast_627_inst_ack_0 : boolean;
  signal type_cast_641_inst_req_1 : boolean;
  signal type_cast_623_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_549_inst_req_0 : boolean;
  signal addr_of_1195_final_reg_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_287_inst_req_1 : boolean;
  signal type_cast_291_inst_req_0 : boolean;
  signal type_cast_291_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_287_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_273_inst_req_0 : boolean;
  signal type_cast_695_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_273_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_587_inst_req_1 : boolean;
  signal type_cast_609_inst_ack_0 : boolean;
  signal type_cast_566_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_287_inst_req_0 : boolean;
  signal type_cast_609_inst_req_0 : boolean;
  signal call_stmt_1072_call_ack_0 : boolean;
  signal phi_stmt_712_req_1 : boolean;
  signal type_cast_745_inst_req_1 : boolean;
  signal type_cast_609_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_299_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_299_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_312_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_312_inst_ack_1 : boolean;
  signal call_stmt_1072_call_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_574_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_741_inst_req_0 : boolean;
  signal type_cast_566_inst_ack_1 : boolean;
  signal type_cast_303_inst_req_1 : boolean;
  signal type_cast_695_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_299_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_312_inst_ack_0 : boolean;
  signal type_cast_316_inst_req_0 : boolean;
  signal type_cast_316_inst_ack_0 : boolean;
  signal type_cast_316_inst_req_1 : boolean;
  signal type_cast_316_inst_ack_1 : boolean;
  signal type_cast_303_inst_ack_1 : boolean;
  signal type_cast_641_inst_ack_1 : boolean;
  signal ptr_deref_1219_store_0_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_549_inst_ack_0 : boolean;
  signal type_cast_278_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_273_inst_ack_1 : boolean;
  signal array_obj_ref_724_index_offset_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_312_inst_req_0 : boolean;
  signal type_cast_623_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_587_inst_ack_1 : boolean;
  signal type_cast_541_inst_req_0 : boolean;
  signal type_cast_623_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_549_inst_req_1 : boolean;
  signal type_cast_278_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_549_inst_ack_1 : boolean;
  signal addr_of_725_final_reg_req_0 : boolean;
  signal type_cast_578_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_574_inst_req_1 : boolean;
  signal type_cast_645_inst_req_0 : boolean;
  signal type_cast_645_inst_req_1 : boolean;
  signal type_cast_278_inst_ack_0 : boolean;
  signal type_cast_645_inst_ack_0 : boolean;
  signal type_cast_541_inst_req_1 : boolean;
  signal if_stmt_668_branch_req_0 : boolean;
  signal type_cast_278_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_537_inst_ack_1 : boolean;
  signal type_cast_627_inst_req_1 : boolean;
  signal type_cast_745_inst_ack_1 : boolean;
  signal type_cast_541_inst_ack_1 : boolean;
  signal type_cast_627_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_741_inst_ack_1 : boolean;
  signal type_cast_1235_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_741_inst_ack_0 : boolean;
  signal array_obj_ref_1215_index_offset_req_1 : boolean;
  signal array_obj_ref_1215_index_offset_req_0 : boolean;
  signal type_cast_732_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_741_inst_req_1 : boolean;
  signal array_obj_ref_724_index_offset_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_324_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_324_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_562_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_324_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_324_inst_ack_1 : boolean;
  signal type_cast_745_inst_ack_0 : boolean;
  signal type_cast_605_inst_ack_0 : boolean;
  signal type_cast_605_inst_req_0 : boolean;
  signal type_cast_328_inst_req_0 : boolean;
  signal type_cast_328_inst_ack_0 : boolean;
  signal array_obj_ref_1215_index_offset_ack_0 : boolean;
  signal type_cast_328_inst_req_1 : boolean;
  signal type_cast_328_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_562_inst_req_1 : boolean;
  signal addr_of_1195_final_reg_req_1 : boolean;
  signal array_obj_ref_724_index_offset_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_337_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_337_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_337_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_337_inst_ack_1 : boolean;
  signal type_cast_745_inst_req_0 : boolean;
  signal type_cast_601_inst_ack_1 : boolean;
  signal type_cast_601_inst_req_1 : boolean;
  signal type_cast_341_inst_req_0 : boolean;
  signal type_cast_341_inst_ack_0 : boolean;
  signal type_cast_341_inst_req_1 : boolean;
  signal type_cast_341_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_562_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_562_inst_req_0 : boolean;
  signal array_obj_ref_724_index_offset_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_349_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_349_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_349_inst_req_1 : boolean;
  signal call_stmt_1290_call_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_349_inst_ack_1 : boolean;
  signal ptr_deref_1199_load_0_ack_0 : boolean;
  signal type_cast_601_inst_ack_0 : boolean;
  signal type_cast_601_inst_req_0 : boolean;
  signal type_cast_353_inst_req_0 : boolean;
  signal if_stmt_668_branch_ack_0 : boolean;
  signal type_cast_353_inst_ack_0 : boolean;
  signal type_cast_353_inst_req_1 : boolean;
  signal type_cast_353_inst_ack_1 : boolean;
  signal addr_of_1195_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_362_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_362_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_362_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_362_inst_ack_1 : boolean;
  signal type_cast_732_inst_ack_1 : boolean;
  signal type_cast_732_inst_req_1 : boolean;
  signal type_cast_366_inst_req_0 : boolean;
  signal type_cast_366_inst_ack_0 : boolean;
  signal type_cast_366_inst_req_1 : boolean;
  signal type_cast_366_inst_ack_1 : boolean;
  signal type_cast_553_inst_ack_1 : boolean;
  signal type_cast_553_inst_req_1 : boolean;
  signal type_cast_591_inst_ack_1 : boolean;
  signal type_cast_591_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_374_inst_req_0 : boolean;
  signal if_stmt_668_branch_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_374_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_374_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_374_inst_ack_1 : boolean;
  signal type_cast_732_inst_ack_0 : boolean;
  signal type_cast_591_inst_ack_0 : boolean;
  signal type_cast_591_inst_req_0 : boolean;
  signal type_cast_378_inst_req_0 : boolean;
  signal type_cast_378_inst_ack_0 : boolean;
  signal type_cast_378_inst_req_1 : boolean;
  signal type_cast_378_inst_ack_1 : boolean;
  signal type_cast_553_inst_ack_0 : boolean;
  signal type_cast_553_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_387_inst_req_0 : boolean;
  signal call_stmt_1290_call_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_387_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_387_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_387_inst_ack_1 : boolean;
  signal call_stmt_1072_call_req_1 : boolean;
  signal type_cast_391_inst_req_0 : boolean;
  signal type_cast_391_inst_ack_0 : boolean;
  signal type_cast_391_inst_req_1 : boolean;
  signal type_cast_391_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_399_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_399_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_399_inst_req_1 : boolean;
  signal call_stmt_1290_call_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_399_inst_ack_1 : boolean;
  signal type_cast_403_inst_req_0 : boolean;
  signal type_cast_403_inst_ack_0 : boolean;
  signal type_cast_403_inst_req_1 : boolean;
  signal type_cast_403_inst_ack_1 : boolean;
  signal addr_of_1216_final_reg_req_0 : boolean;
  signal addr_of_1216_final_reg_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_412_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_412_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_412_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_412_inst_ack_1 : boolean;
  signal addr_of_1216_final_reg_req_1 : boolean;
  signal addr_of_1216_final_reg_ack_1 : boolean;
  signal type_cast_416_inst_req_0 : boolean;
  signal type_cast_416_inst_ack_0 : boolean;
  signal type_cast_416_inst_req_1 : boolean;
  signal type_cast_416_inst_ack_1 : boolean;
  signal type_cast_1235_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_424_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_424_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_424_inst_req_1 : boolean;
  signal call_stmt_1290_call_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_424_inst_ack_1 : boolean;
  signal phi_stmt_950_req_1 : boolean;
  signal type_cast_428_inst_req_0 : boolean;
  signal type_cast_428_inst_ack_0 : boolean;
  signal type_cast_428_inst_req_1 : boolean;
  signal type_cast_428_inst_ack_1 : boolean;
  signal call_stmt_1072_call_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_437_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_437_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_437_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_437_inst_ack_1 : boolean;
  signal type_cast_1235_inst_ack_0 : boolean;
  signal type_cast_441_inst_req_0 : boolean;
  signal type_cast_441_inst_ack_0 : boolean;
  signal type_cast_441_inst_req_1 : boolean;
  signal type_cast_441_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_449_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_449_inst_ack_0 : boolean;
  signal type_cast_956_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_449_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_449_inst_ack_1 : boolean;
  signal type_cast_453_inst_req_0 : boolean;
  signal type_cast_453_inst_ack_0 : boolean;
  signal type_cast_453_inst_req_1 : boolean;
  signal type_cast_453_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_462_inst_req_0 : boolean;
  signal type_cast_1294_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_462_inst_ack_0 : boolean;
  signal type_cast_1294_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_462_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_462_inst_ack_1 : boolean;
  signal phi_stmt_950_req_0 : boolean;
  signal type_cast_466_inst_req_0 : boolean;
  signal type_cast_466_inst_ack_0 : boolean;
  signal type_cast_466_inst_req_1 : boolean;
  signal type_cast_466_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_474_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_474_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_474_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_474_inst_ack_1 : boolean;
  signal type_cast_478_inst_req_0 : boolean;
  signal type_cast_478_inst_ack_0 : boolean;
  signal type_cast_478_inst_req_1 : boolean;
  signal type_cast_478_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_487_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_487_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_487_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_487_inst_ack_1 : boolean;
  signal type_cast_491_inst_req_0 : boolean;
  signal type_cast_491_inst_ack_0 : boolean;
  signal type_cast_491_inst_req_1 : boolean;
  signal type_cast_491_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_499_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_499_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_499_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_499_inst_ack_1 : boolean;
  signal type_cast_503_inst_req_0 : boolean;
  signal type_cast_503_inst_ack_0 : boolean;
  signal type_cast_503_inst_req_1 : boolean;
  signal type_cast_503_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_512_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_512_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_512_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_512_inst_ack_1 : boolean;
  signal type_cast_516_inst_req_0 : boolean;
  signal type_cast_516_inst_ack_0 : boolean;
  signal type_cast_516_inst_req_1 : boolean;
  signal type_cast_516_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_524_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_524_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_524_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_524_inst_ack_1 : boolean;
  signal type_cast_528_inst_req_0 : boolean;
  signal type_cast_528_inst_ack_0 : boolean;
  signal type_cast_528_inst_req_1 : boolean;
  signal type_cast_528_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_537_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_537_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_759_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_759_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_759_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_759_inst_ack_1 : boolean;
  signal type_cast_718_inst_ack_1 : boolean;
  signal type_cast_763_inst_req_0 : boolean;
  signal type_cast_763_inst_ack_0 : boolean;
  signal type_cast_763_inst_req_1 : boolean;
  signal type_cast_1286_inst_ack_1 : boolean;
  signal type_cast_763_inst_ack_1 : boolean;
  signal phi_stmt_950_ack_0 : boolean;
  signal type_cast_718_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_777_inst_req_0 : boolean;
  signal type_cast_1286_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_777_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_777_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_777_inst_ack_1 : boolean;
  signal type_cast_956_inst_ack_1 : boolean;
  signal type_cast_781_inst_req_0 : boolean;
  signal type_cast_781_inst_ack_0 : boolean;
  signal type_cast_781_inst_req_1 : boolean;
  signal type_cast_1286_inst_ack_0 : boolean;
  signal type_cast_781_inst_ack_1 : boolean;
  signal array_obj_ref_1194_index_offset_ack_1 : boolean;
  signal array_obj_ref_1194_index_offset_req_1 : boolean;
  signal type_cast_718_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_795_inst_req_0 : boolean;
  signal type_cast_1286_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_795_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_795_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_795_inst_ack_1 : boolean;
  signal type_cast_799_inst_req_0 : boolean;
  signal type_cast_799_inst_ack_0 : boolean;
  signal type_cast_799_inst_req_1 : boolean;
  signal type_cast_799_inst_ack_1 : boolean;
  signal type_cast_718_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_813_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_813_inst_ack_0 : boolean;
  signal array_obj_ref_1194_index_offset_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_813_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_813_inst_ack_1 : boolean;
  signal type_cast_956_inst_req_1 : boolean;
  signal call_stmt_1306_call_ack_1 : boolean;
  signal type_cast_817_inst_req_0 : boolean;
  signal type_cast_817_inst_ack_0 : boolean;
  signal type_cast_817_inst_req_1 : boolean;
  signal type_cast_817_inst_ack_1 : boolean;
  signal call_stmt_1306_call_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_831_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_831_inst_ack_0 : boolean;
  signal array_obj_ref_1194_index_offset_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_831_inst_req_1 : boolean;
  signal if_stmt_1275_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_831_inst_ack_1 : boolean;
  signal type_cast_835_inst_req_0 : boolean;
  signal type_cast_835_inst_ack_0 : boolean;
  signal type_cast_835_inst_req_1 : boolean;
  signal type_cast_835_inst_ack_1 : boolean;
  signal call_stmt_1306_call_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_849_inst_req_0 : boolean;
  signal if_stmt_1275_branch_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_849_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_849_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_849_inst_ack_1 : boolean;
  signal call_stmt_1306_call_req_0 : boolean;
  signal type_cast_853_inst_req_0 : boolean;
  signal type_cast_853_inst_ack_0 : boolean;
  signal type_cast_853_inst_req_1 : boolean;
  signal if_stmt_1275_branch_req_0 : boolean;
  signal type_cast_853_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1301_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1301_inst_req_1 : boolean;
  signal ptr_deref_1199_load_0_req_0 : boolean;
  signal ptr_deref_861_store_0_req_0 : boolean;
  signal ptr_deref_861_store_0_ack_0 : boolean;
  signal ptr_deref_1219_store_0_ack_0 : boolean;
  signal ptr_deref_861_store_0_req_1 : boolean;
  signal ptr_deref_861_store_0_ack_1 : boolean;
  signal ptr_deref_1219_store_0_req_0 : boolean;
  signal if_stmt_875_branch_req_0 : boolean;
  signal type_cast_1203_inst_ack_1 : boolean;
  signal if_stmt_875_branch_ack_1 : boolean;
  signal if_stmt_875_branch_ack_0 : boolean;
  signal if_stmt_891_branch_req_0 : boolean;
  signal type_cast_1203_inst_req_1 : boolean;
  signal type_cast_1182_inst_ack_1 : boolean;
  signal type_cast_1182_inst_req_1 : boolean;
  signal if_stmt_891_branch_ack_1 : boolean;
  signal if_stmt_891_branch_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1301_inst_ack_0 : boolean;
  signal type_cast_933_inst_req_0 : boolean;
  signal type_cast_1256_inst_ack_1 : boolean;
  signal type_cast_933_inst_ack_0 : boolean;
  signal type_cast_933_inst_req_1 : boolean;
  signal type_cast_1256_inst_req_1 : boolean;
  signal type_cast_933_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1301_inst_req_0 : boolean;
  signal call_stmt_959_call_req_0 : boolean;
  signal call_stmt_959_call_ack_0 : boolean;
  signal call_stmt_959_call_req_1 : boolean;
  signal call_stmt_959_call_ack_1 : boolean;
  signal type_cast_1182_inst_ack_0 : boolean;
  signal if_stmt_971_branch_req_0 : boolean;
  signal type_cast_1182_inst_req_0 : boolean;
  signal if_stmt_971_branch_ack_1 : boolean;
  signal if_stmt_971_branch_ack_0 : boolean;
  signal type_cast_1256_inst_ack_0 : boolean;
  signal if_stmt_987_branch_req_0 : boolean;
  signal type_cast_1203_inst_ack_0 : boolean;
  signal if_stmt_987_branch_ack_1 : boolean;
  signal if_stmt_987_branch_ack_0 : boolean;
  signal phi_stmt_712_ack_0 : boolean;
  signal type_cast_1014_inst_req_0 : boolean;
  signal type_cast_1256_inst_req_0 : boolean;
  signal type_cast_1014_inst_ack_0 : boolean;
  signal type_cast_1014_inst_req_1 : boolean;
  signal type_cast_1014_inst_ack_1 : boolean;
  signal phi_stmt_712_req_0 : boolean;
  signal type_cast_1203_inst_req_0 : boolean;
  signal type_cast_1294_inst_ack_1 : boolean;
  signal type_cast_956_inst_ack_0 : boolean;
  signal array_obj_ref_1043_index_offset_req_0 : boolean;
  signal array_obj_ref_1043_index_offset_ack_0 : boolean;
  signal array_obj_ref_1043_index_offset_req_1 : boolean;
  signal array_obj_ref_1043_index_offset_ack_1 : boolean;
  signal addr_of_1044_final_reg_req_0 : boolean;
  signal addr_of_1044_final_reg_ack_0 : boolean;
  signal addr_of_1044_final_reg_req_1 : boolean;
  signal type_cast_1235_inst_ack_1 : boolean;
  signal addr_of_1044_final_reg_ack_1 : boolean;
  signal type_cast_1294_inst_req_1 : boolean;
  signal ptr_deref_1199_load_0_ack_1 : boolean;
  signal ptr_deref_1199_load_0_req_1 : boolean;
  signal ptr_deref_1047_store_0_req_0 : boolean;
  signal ptr_deref_1047_store_0_ack_0 : boolean;
  signal ptr_deref_1047_store_0_req_1 : boolean;
  signal ptr_deref_1047_store_0_ack_1 : boolean;
  signal if_stmt_1062_branch_req_0 : boolean;
  signal if_stmt_1062_branch_ack_1 : boolean;
  signal if_stmt_1062_branch_ack_0 : boolean;
  signal phi_stmt_1031_req_0 : boolean;
  signal type_cast_1037_inst_req_0 : boolean;
  signal type_cast_1037_inst_ack_0 : boolean;
  signal type_cast_1037_inst_req_1 : boolean;
  signal type_cast_1037_inst_ack_1 : boolean;
  signal phi_stmt_1031_req_1 : boolean;
  signal phi_stmt_1031_ack_0 : boolean;
  signal phi_stmt_1098_req_0 : boolean;
  signal phi_stmt_1105_req_0 : boolean;
  signal phi_stmt_1112_req_0 : boolean;
  signal type_cast_1104_inst_req_0 : boolean;
  signal type_cast_1104_inst_ack_0 : boolean;
  signal type_cast_1104_inst_req_1 : boolean;
  signal type_cast_1104_inst_ack_1 : boolean;
  signal phi_stmt_1098_req_1 : boolean;
  signal type_cast_1111_inst_req_0 : boolean;
  signal type_cast_1111_inst_ack_0 : boolean;
  signal type_cast_1111_inst_req_1 : boolean;
  signal type_cast_1111_inst_ack_1 : boolean;
  signal phi_stmt_1105_req_1 : boolean;
  signal type_cast_1118_inst_req_0 : boolean;
  signal type_cast_1118_inst_ack_0 : boolean;
  signal type_cast_1118_inst_req_1 : boolean;
  signal type_cast_1118_inst_ack_1 : boolean;
  signal phi_stmt_1112_req_1 : boolean;
  signal phi_stmt_1098_ack_0 : boolean;
  signal phi_stmt_1105_ack_0 : boolean;
  signal phi_stmt_1112_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_814_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_814_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_814_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_814_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_814: Block -- control-path 
    signal convTranspose_CP_814_elements: BooleanArray(263 downto 0);
    -- 
  begin -- 
    convTranspose_CP_814_elements(0) <= convTranspose_CP_814_start;
    convTranspose_CP_814_symbol <= convTranspose_CP_814_elements(223);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	72 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	64 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	68 
    -- CP-element group 0: 	80 
    -- CP-element group 0: 	96 
    -- CP-element group 0: 	88 
    -- CP-element group 0: 	100 
    -- CP-element group 0: 	76 
    -- CP-element group 0: 	84 
    -- CP-element group 0: 	104 
    -- CP-element group 0: 	92 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0:  members (86) 
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_566_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597__entry__
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_541_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_578_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/branch_block_stmt_271__entry__
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_553_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_316_update_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_578_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_566_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_291_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_273_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_273_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_273_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_303_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_303_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_303_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_291_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_566_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_316_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_316_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_291_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_278_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_278_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_541_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_541_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_278_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_578_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_328_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_328_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_328_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_341_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_341_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_341_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_353_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_353_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_353_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_366_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_366_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_366_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_553_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_591_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_553_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_591_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_378_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_378_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_378_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_591_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_391_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_391_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_391_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_403_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_403_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_403_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_416_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_416_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_416_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_428_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_428_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_428_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_441_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_441_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_441_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_453_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_453_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_453_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_466_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_466_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_466_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_478_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_478_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_478_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_491_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_491_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_491_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_503_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_503_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_503_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_516_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_516_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_516_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_528_update_start_
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_528_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_528_Update/cr
      -- 
    cr_1571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_566_inst_req_1); -- 
    cr_1599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_578_inst_req_1); -- 
    cr_955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_291_inst_req_1); -- 
    rr_908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => RPIPE_ConvTranspose_input_pipe_273_inst_req_0); -- 
    cr_983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_303_inst_req_1); -- 
    cr_1011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_316_inst_req_1); -- 
    cr_927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_278_inst_req_1); -- 
    cr_1515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_541_inst_req_1); -- 
    cr_1039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_328_inst_req_1); -- 
    cr_1067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_341_inst_req_1); -- 
    cr_1095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_353_inst_req_1); -- 
    cr_1123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_366_inst_req_1); -- 
    cr_1543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_553_inst_req_1); -- 
    cr_1627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_591_inst_req_1); -- 
    cr_1151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_378_inst_req_1); -- 
    cr_1179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_391_inst_req_1); -- 
    cr_1207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_403_inst_req_1); -- 
    cr_1235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_416_inst_req_1); -- 
    cr_1263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_428_inst_req_1); -- 
    cr_1291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_441_inst_req_1); -- 
    cr_1319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_453_inst_req_1); -- 
    cr_1347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_466_inst_req_1); -- 
    cr_1375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_478_inst_req_1); -- 
    cr_1403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_491_inst_req_1); -- 
    cr_1431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_503_inst_req_1); -- 
    cr_1459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_516_inst_req_1); -- 
    cr_1487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(0), ack => type_cast_528_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_273_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_273_update_start_
      -- CP-element group 1: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_273_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_273_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_273_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_273_Update/$entry
      -- 
    ra_909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_273_inst_ack_0, ack => convTranspose_CP_814_elements(1)); -- 
    cr_913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(1), ack => RPIPE_ConvTranspose_input_pipe_273_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_287_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_273_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_287_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_278_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_287_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_273_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_273_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_278_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_278_Sample/$entry
      -- 
    ca_914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_273_inst_ack_1, ack => convTranspose_CP_814_elements(2)); -- 
    rr_922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(2), ack => type_cast_278_inst_req_0); -- 
    rr_936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(2), ack => RPIPE_ConvTranspose_input_pipe_287_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_278_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_278_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_278_Sample/$exit
      -- 
    ra_923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_278_inst_ack_0, ack => convTranspose_CP_814_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	105 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_278_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_278_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_278_update_completed_
      -- 
    ca_928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_278_inst_ack_1, ack => convTranspose_CP_814_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_287_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_287_Update/cr
      -- CP-element group 5: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_287_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_287_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_287_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_287_update_start_
      -- 
    ra_937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_287_inst_ack_0, ack => convTranspose_CP_814_elements(5)); -- 
    cr_941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(5), ack => RPIPE_ConvTranspose_input_pipe_287_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_287_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_291_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_287_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_287_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_299_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_299_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_291_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_299_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_291_Sample/$entry
      -- 
    ca_942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_287_inst_ack_1, ack => convTranspose_CP_814_elements(6)); -- 
    rr_950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(6), ack => type_cast_291_inst_req_0); -- 
    rr_964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(6), ack => RPIPE_ConvTranspose_input_pipe_299_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_291_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_291_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_291_sample_completed_
      -- 
    ra_951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_291_inst_ack_0, ack => convTranspose_CP_814_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	105 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_291_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_291_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_291_update_completed_
      -- 
    ca_956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_291_inst_ack_1, ack => convTranspose_CP_814_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_299_Update/cr
      -- CP-element group 9: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_299_update_start_
      -- CP-element group 9: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_299_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_299_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_299_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_299_Update/$entry
      -- 
    ra_965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_299_inst_ack_0, ack => convTranspose_CP_814_elements(9)); -- 
    cr_969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(9), ack => RPIPE_ConvTranspose_input_pipe_299_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_303_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_299_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_303_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_299_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_303_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_299_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_312_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_312_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_312_Sample/rr
      -- 
    ca_970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_299_inst_ack_1, ack => convTranspose_CP_814_elements(10)); -- 
    rr_978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(10), ack => type_cast_303_inst_req_0); -- 
    rr_992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(10), ack => RPIPE_ConvTranspose_input_pipe_312_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_303_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_303_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_303_Sample/$exit
      -- 
    ra_979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_303_inst_ack_0, ack => convTranspose_CP_814_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	105 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_303_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_303_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_303_Update/ca
      -- 
    ca_984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_303_inst_ack_1, ack => convTranspose_CP_814_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_312_Update/cr
      -- CP-element group 13: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_312_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_312_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_312_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_312_update_start_
      -- CP-element group 13: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_312_Sample/$exit
      -- 
    ra_993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_312_inst_ack_0, ack => convTranspose_CP_814_elements(13)); -- 
    cr_997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(13), ack => RPIPE_ConvTranspose_input_pipe_312_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_312_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_316_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_312_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_316_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_316_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_312_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_324_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_324_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_324_Sample/rr
      -- 
    ca_998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_312_inst_ack_1, ack => convTranspose_CP_814_elements(14)); -- 
    rr_1006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(14), ack => type_cast_316_inst_req_0); -- 
    rr_1020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(14), ack => RPIPE_ConvTranspose_input_pipe_324_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_316_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_316_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_316_Sample/ra
      -- 
    ra_1007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_316_inst_ack_0, ack => convTranspose_CP_814_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	105 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_316_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_316_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_316_Update/ca
      -- 
    ca_1012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_316_inst_ack_1, ack => convTranspose_CP_814_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_324_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_324_update_start_
      -- CP-element group 17: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_324_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_324_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_324_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_324_Update/cr
      -- 
    ra_1021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_324_inst_ack_0, ack => convTranspose_CP_814_elements(17)); -- 
    cr_1025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(17), ack => RPIPE_ConvTranspose_input_pipe_324_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_324_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_324_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_324_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_328_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_328_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_328_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_337_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_337_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_337_Sample/rr
      -- 
    ca_1026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_324_inst_ack_1, ack => convTranspose_CP_814_elements(18)); -- 
    rr_1034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(18), ack => type_cast_328_inst_req_0); -- 
    rr_1048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(18), ack => RPIPE_ConvTranspose_input_pipe_337_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_328_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_328_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_328_Sample/ra
      -- 
    ra_1035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_328_inst_ack_0, ack => convTranspose_CP_814_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	105 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_328_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_328_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_328_Update/ca
      -- 
    ca_1040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_328_inst_ack_1, ack => convTranspose_CP_814_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_337_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_337_update_start_
      -- CP-element group 21: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_337_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_337_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_337_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_337_Update/cr
      -- 
    ra_1049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_337_inst_ack_0, ack => convTranspose_CP_814_elements(21)); -- 
    cr_1053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(21), ack => RPIPE_ConvTranspose_input_pipe_337_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_337_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_337_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_337_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_341_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_341_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_341_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_349_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_349_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_349_Sample/rr
      -- 
    ca_1054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_337_inst_ack_1, ack => convTranspose_CP_814_elements(22)); -- 
    rr_1062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(22), ack => type_cast_341_inst_req_0); -- 
    rr_1076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(22), ack => RPIPE_ConvTranspose_input_pipe_349_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_341_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_341_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_341_Sample/ra
      -- 
    ra_1063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_341_inst_ack_0, ack => convTranspose_CP_814_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	105 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_341_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_341_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_341_Update/ca
      -- 
    ca_1068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_341_inst_ack_1, ack => convTranspose_CP_814_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_349_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_349_update_start_
      -- CP-element group 25: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_349_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_349_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_349_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_349_Update/cr
      -- 
    ra_1077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_349_inst_ack_0, ack => convTranspose_CP_814_elements(25)); -- 
    cr_1081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(25), ack => RPIPE_ConvTranspose_input_pipe_349_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_349_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_349_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_349_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_353_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_353_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_353_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_362_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_362_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_362_Sample/rr
      -- 
    ca_1082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_349_inst_ack_1, ack => convTranspose_CP_814_elements(26)); -- 
    rr_1090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(26), ack => type_cast_353_inst_req_0); -- 
    rr_1104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(26), ack => RPIPE_ConvTranspose_input_pipe_362_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_353_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_353_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_353_Sample/ra
      -- 
    ra_1091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_353_inst_ack_0, ack => convTranspose_CP_814_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	105 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_353_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_353_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_353_Update/ca
      -- 
    ca_1096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_353_inst_ack_1, ack => convTranspose_CP_814_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_362_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_362_update_start_
      -- CP-element group 29: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_362_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_362_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_362_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_362_Update/cr
      -- 
    ra_1105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_362_inst_ack_0, ack => convTranspose_CP_814_elements(29)); -- 
    cr_1109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(29), ack => RPIPE_ConvTranspose_input_pipe_362_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	33 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_362_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_362_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_362_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_366_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_366_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_366_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_374_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_374_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_374_Sample/rr
      -- 
    ca_1110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_362_inst_ack_1, ack => convTranspose_CP_814_elements(30)); -- 
    rr_1132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(30), ack => RPIPE_ConvTranspose_input_pipe_374_inst_req_0); -- 
    rr_1118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(30), ack => type_cast_366_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_366_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_366_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_366_Sample/ra
      -- 
    ra_1119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_366_inst_ack_0, ack => convTranspose_CP_814_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	105 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_366_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_366_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_366_Update/ca
      -- 
    ca_1124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_366_inst_ack_1, ack => convTranspose_CP_814_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_374_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_374_update_start_
      -- CP-element group 33: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_374_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_374_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_374_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_374_Update/cr
      -- 
    ra_1133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_374_inst_ack_0, ack => convTranspose_CP_814_elements(33)); -- 
    cr_1137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(33), ack => RPIPE_ConvTranspose_input_pipe_374_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_374_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_374_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_374_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_378_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_378_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_378_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_387_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_387_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_387_Sample/rr
      -- 
    ca_1138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_374_inst_ack_1, ack => convTranspose_CP_814_elements(34)); -- 
    rr_1160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(34), ack => RPIPE_ConvTranspose_input_pipe_387_inst_req_0); -- 
    rr_1146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(34), ack => type_cast_378_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_378_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_378_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_378_Sample/ra
      -- 
    ra_1147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_378_inst_ack_0, ack => convTranspose_CP_814_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	105 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_378_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_378_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_378_Update/ca
      -- 
    ca_1152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_378_inst_ack_1, ack => convTranspose_CP_814_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_387_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_387_update_start_
      -- CP-element group 37: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_387_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_387_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_387_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_387_Update/cr
      -- 
    ra_1161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_387_inst_ack_0, ack => convTranspose_CP_814_elements(37)); -- 
    cr_1165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(37), ack => RPIPE_ConvTranspose_input_pipe_387_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_387_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_387_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_387_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_391_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_391_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_391_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_399_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_399_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_399_Sample/rr
      -- 
    ca_1166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_387_inst_ack_1, ack => convTranspose_CP_814_elements(38)); -- 
    rr_1174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(38), ack => type_cast_391_inst_req_0); -- 
    rr_1188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(38), ack => RPIPE_ConvTranspose_input_pipe_399_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_391_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_391_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_391_Sample/ra
      -- 
    ra_1175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_391_inst_ack_0, ack => convTranspose_CP_814_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	105 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_391_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_391_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_391_Update/ca
      -- 
    ca_1180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_391_inst_ack_1, ack => convTranspose_CP_814_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_399_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_399_update_start_
      -- CP-element group 41: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_399_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_399_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_399_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_399_Update/cr
      -- 
    ra_1189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_399_inst_ack_0, ack => convTranspose_CP_814_elements(41)); -- 
    cr_1193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(41), ack => RPIPE_ConvTranspose_input_pipe_399_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	45 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_399_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_399_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_399_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_403_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_403_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_403_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_412_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_412_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_412_Sample/rr
      -- 
    ca_1194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_399_inst_ack_1, ack => convTranspose_CP_814_elements(42)); -- 
    rr_1202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(42), ack => type_cast_403_inst_req_0); -- 
    rr_1216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(42), ack => RPIPE_ConvTranspose_input_pipe_412_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_403_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_403_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_403_Sample/ra
      -- 
    ra_1203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_403_inst_ack_0, ack => convTranspose_CP_814_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	105 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_403_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_403_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_403_Update/ca
      -- 
    ca_1208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_403_inst_ack_1, ack => convTranspose_CP_814_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_412_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_412_update_start_
      -- CP-element group 45: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_412_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_412_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_412_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_412_Update/cr
      -- 
    ra_1217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_412_inst_ack_0, ack => convTranspose_CP_814_elements(45)); -- 
    cr_1221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(45), ack => RPIPE_ConvTranspose_input_pipe_412_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	49 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_412_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_412_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_412_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_416_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_416_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_416_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_424_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_424_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_424_Sample/rr
      -- 
    ca_1222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_412_inst_ack_1, ack => convTranspose_CP_814_elements(46)); -- 
    rr_1230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(46), ack => type_cast_416_inst_req_0); -- 
    rr_1244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(46), ack => RPIPE_ConvTranspose_input_pipe_424_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_416_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_416_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_416_Sample/ra
      -- 
    ra_1231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_416_inst_ack_0, ack => convTranspose_CP_814_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	105 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_416_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_416_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_416_Update/ca
      -- 
    ca_1236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_416_inst_ack_1, ack => convTranspose_CP_814_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_424_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_424_update_start_
      -- CP-element group 49: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_424_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_424_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_424_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_424_Update/cr
      -- 
    ra_1245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_424_inst_ack_0, ack => convTranspose_CP_814_elements(49)); -- 
    cr_1249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(49), ack => RPIPE_ConvTranspose_input_pipe_424_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_424_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_424_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_424_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_428_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_428_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_428_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_437_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_437_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_437_Sample/rr
      -- 
    ca_1250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_424_inst_ack_1, ack => convTranspose_CP_814_elements(50)); -- 
    rr_1258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(50), ack => type_cast_428_inst_req_0); -- 
    rr_1272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(50), ack => RPIPE_ConvTranspose_input_pipe_437_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_428_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_428_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_428_Sample/ra
      -- 
    ra_1259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_428_inst_ack_0, ack => convTranspose_CP_814_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	105 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_428_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_428_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_428_Update/ca
      -- 
    ca_1264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_428_inst_ack_1, ack => convTranspose_CP_814_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_437_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_437_update_start_
      -- CP-element group 53: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_437_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_437_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_437_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_437_Update/cr
      -- 
    ra_1273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_437_inst_ack_0, ack => convTranspose_CP_814_elements(53)); -- 
    cr_1277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(53), ack => RPIPE_ConvTranspose_input_pipe_437_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	57 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_437_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_437_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_437_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_441_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_441_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_441_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_449_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_449_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_449_Sample/rr
      -- 
    ca_1278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_437_inst_ack_1, ack => convTranspose_CP_814_elements(54)); -- 
    rr_1286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(54), ack => type_cast_441_inst_req_0); -- 
    rr_1300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(54), ack => RPIPE_ConvTranspose_input_pipe_449_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_441_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_441_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_441_Sample/ra
      -- 
    ra_1287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_441_inst_ack_0, ack => convTranspose_CP_814_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	105 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_441_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_441_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_441_Update/ca
      -- 
    ca_1292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_441_inst_ack_1, ack => convTranspose_CP_814_elements(56)); -- 
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	54 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_449_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_449_update_start_
      -- CP-element group 57: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_449_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_449_Sample/ra
      -- CP-element group 57: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_449_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_449_Update/cr
      -- 
    ra_1301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_449_inst_ack_0, ack => convTranspose_CP_814_elements(57)); -- 
    cr_1305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(57), ack => RPIPE_ConvTranspose_input_pipe_449_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	61 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_449_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_449_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_449_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_453_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_453_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_453_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_462_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_462_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_462_Sample/rr
      -- 
    ca_1306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_449_inst_ack_1, ack => convTranspose_CP_814_elements(58)); -- 
    rr_1328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(58), ack => RPIPE_ConvTranspose_input_pipe_462_inst_req_0); -- 
    rr_1314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(58), ack => type_cast_453_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_453_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_453_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_453_Sample/ra
      -- 
    ra_1315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_453_inst_ack_0, ack => convTranspose_CP_814_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	105 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_453_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_453_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_453_Update/ca
      -- 
    ca_1320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_453_inst_ack_1, ack => convTranspose_CP_814_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	58 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_462_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_462_update_start_
      -- CP-element group 61: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_462_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_462_Sample/ra
      -- CP-element group 61: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_462_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_462_Update/cr
      -- 
    ra_1329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_462_inst_ack_0, ack => convTranspose_CP_814_elements(61)); -- 
    cr_1333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(61), ack => RPIPE_ConvTranspose_input_pipe_462_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	65 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (9) 
      -- CP-element group 62: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_462_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_462_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_462_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_466_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_466_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_466_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_474_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_474_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_474_Sample/rr
      -- 
    ca_1334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_462_inst_ack_1, ack => convTranspose_CP_814_elements(62)); -- 
    rr_1342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(62), ack => type_cast_466_inst_req_0); -- 
    rr_1356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(62), ack => RPIPE_ConvTranspose_input_pipe_474_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_466_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_466_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_466_Sample/ra
      -- 
    ra_1343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_466_inst_ack_0, ack => convTranspose_CP_814_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	0 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	105 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_466_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_466_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_466_Update/ca
      -- 
    ca_1348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_466_inst_ack_1, ack => convTranspose_CP_814_elements(64)); -- 
    -- CP-element group 65:  transition  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	62 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (6) 
      -- CP-element group 65: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_474_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_474_update_start_
      -- CP-element group 65: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_474_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_474_Sample/ra
      -- CP-element group 65: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_474_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_474_Update/cr
      -- 
    ra_1357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_474_inst_ack_0, ack => convTranspose_CP_814_elements(65)); -- 
    cr_1361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(65), ack => RPIPE_ConvTranspose_input_pipe_474_inst_req_1); -- 
    -- CP-element group 66:  fork  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	69 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (9) 
      -- CP-element group 66: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_474_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_474_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_474_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_478_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_478_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_478_Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_487_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_487_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_487_Sample/rr
      -- 
    ca_1362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_474_inst_ack_1, ack => convTranspose_CP_814_elements(66)); -- 
    rr_1370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(66), ack => type_cast_478_inst_req_0); -- 
    rr_1384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(66), ack => RPIPE_ConvTranspose_input_pipe_487_inst_req_0); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_478_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_478_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_478_Sample/ra
      -- 
    ra_1371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_478_inst_ack_0, ack => convTranspose_CP_814_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	0 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	105 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_478_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_478_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_478_Update/ca
      -- 
    ca_1376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_478_inst_ack_1, ack => convTranspose_CP_814_elements(68)); -- 
    -- CP-element group 69:  transition  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	66 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (6) 
      -- CP-element group 69: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_487_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_487_update_start_
      -- CP-element group 69: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_487_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_487_Sample/ra
      -- CP-element group 69: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_487_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_487_Update/cr
      -- 
    ra_1385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_487_inst_ack_0, ack => convTranspose_CP_814_elements(69)); -- 
    cr_1389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(69), ack => RPIPE_ConvTranspose_input_pipe_487_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	73 
    -- CP-element group 70:  members (9) 
      -- CP-element group 70: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_487_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_487_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_487_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_491_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_491_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_491_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_499_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_499_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_499_Sample/rr
      -- 
    ca_1390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_487_inst_ack_1, ack => convTranspose_CP_814_elements(70)); -- 
    rr_1398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(70), ack => type_cast_491_inst_req_0); -- 
    rr_1412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(70), ack => RPIPE_ConvTranspose_input_pipe_499_inst_req_0); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_491_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_491_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_491_Sample/ra
      -- 
    ra_1399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_491_inst_ack_0, ack => convTranspose_CP_814_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	0 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	105 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_491_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_491_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_491_Update/ca
      -- 
    ca_1404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_491_inst_ack_1, ack => convTranspose_CP_814_elements(72)); -- 
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	70 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_499_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_499_update_start_
      -- CP-element group 73: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_499_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_499_Sample/ra
      -- CP-element group 73: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_499_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_499_Update/cr
      -- 
    ra_1413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_499_inst_ack_0, ack => convTranspose_CP_814_elements(73)); -- 
    cr_1417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(73), ack => RPIPE_ConvTranspose_input_pipe_499_inst_req_1); -- 
    -- CP-element group 74:  fork  transition  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	77 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (9) 
      -- CP-element group 74: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_499_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_499_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_499_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_503_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_503_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_503_Sample/rr
      -- CP-element group 74: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_512_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_512_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_512_Sample/rr
      -- 
    ca_1418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_499_inst_ack_1, ack => convTranspose_CP_814_elements(74)); -- 
    rr_1426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(74), ack => type_cast_503_inst_req_0); -- 
    rr_1440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(74), ack => RPIPE_ConvTranspose_input_pipe_512_inst_req_0); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_503_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_503_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_503_Sample/ra
      -- 
    ra_1427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_503_inst_ack_0, ack => convTranspose_CP_814_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	0 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	105 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_503_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_503_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_503_Update/ca
      -- 
    ca_1432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_503_inst_ack_1, ack => convTranspose_CP_814_elements(76)); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	74 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_512_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_512_update_start_
      -- CP-element group 77: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_512_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_512_Sample/ra
      -- CP-element group 77: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_512_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_512_Update/cr
      -- 
    ra_1441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_512_inst_ack_0, ack => convTranspose_CP_814_elements(77)); -- 
    cr_1445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(77), ack => RPIPE_ConvTranspose_input_pipe_512_inst_req_1); -- 
    -- CP-element group 78:  fork  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	81 
    -- CP-element group 78:  members (9) 
      -- CP-element group 78: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_512_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_512_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_512_Update/ca
      -- CP-element group 78: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_516_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_516_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_516_Sample/rr
      -- CP-element group 78: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_524_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_524_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_524_Sample/rr
      -- 
    ca_1446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_512_inst_ack_1, ack => convTranspose_CP_814_elements(78)); -- 
    rr_1454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(78), ack => type_cast_516_inst_req_0); -- 
    rr_1468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(78), ack => RPIPE_ConvTranspose_input_pipe_524_inst_req_0); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_516_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_516_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_516_Sample/ra
      -- 
    ra_1455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_516_inst_ack_0, ack => convTranspose_CP_814_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	0 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	105 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_516_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_516_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_516_Update/ca
      -- 
    ca_1460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_516_inst_ack_1, ack => convTranspose_CP_814_elements(80)); -- 
    -- CP-element group 81:  transition  input  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	78 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (6) 
      -- CP-element group 81: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_524_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_524_update_start_
      -- CP-element group 81: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_524_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_524_Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_524_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_524_Update/cr
      -- 
    ra_1469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_524_inst_ack_0, ack => convTranspose_CP_814_elements(81)); -- 
    cr_1473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(81), ack => RPIPE_ConvTranspose_input_pipe_524_inst_req_1); -- 
    -- CP-element group 82:  fork  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82: 	85 
    -- CP-element group 82:  members (9) 
      -- CP-element group 82: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_524_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_524_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_524_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_528_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_528_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_528_Sample/rr
      -- CP-element group 82: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_537_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_537_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_537_Sample/rr
      -- 
    ca_1474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_524_inst_ack_1, ack => convTranspose_CP_814_elements(82)); -- 
    rr_1482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(82), ack => type_cast_528_inst_req_0); -- 
    rr_1496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(82), ack => RPIPE_ConvTranspose_input_pipe_537_inst_req_0); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_528_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_528_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_528_Sample/ra
      -- 
    ra_1483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_528_inst_ack_0, ack => convTranspose_CP_814_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	0 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	105 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_528_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_528_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_528_Update/ca
      -- 
    ca_1488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_528_inst_ack_1, ack => convTranspose_CP_814_elements(84)); -- 
    -- CP-element group 85:  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	82 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (6) 
      -- CP-element group 85: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_537_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_537_Update/cr
      -- CP-element group 85: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_537_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_537_update_start_
      -- CP-element group 85: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_537_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_537_Sample/ra
      -- 
    ra_1497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_537_inst_ack_0, ack => convTranspose_CP_814_elements(85)); -- 
    cr_1501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(85), ack => RPIPE_ConvTranspose_input_pipe_537_inst_req_1); -- 
    -- CP-element group 86:  fork  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86: 	89 
    -- CP-element group 86:  members (9) 
      -- CP-element group 86: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_549_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_549_Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_541_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_541_Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_537_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_537_Update/ca
      -- CP-element group 86: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_549_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_541_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_537_update_completed_
      -- 
    ca_1502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_537_inst_ack_1, ack => convTranspose_CP_814_elements(86)); -- 
    rr_1510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(86), ack => type_cast_541_inst_req_0); -- 
    rr_1524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(86), ack => RPIPE_ConvTranspose_input_pipe_549_inst_req_0); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_541_Sample/ra
      -- CP-element group 87: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_541_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_541_Sample/$exit
      -- 
    ra_1511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_541_inst_ack_0, ack => convTranspose_CP_814_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	0 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	105 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_541_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_541_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_541_Update/ca
      -- 
    ca_1516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_541_inst_ack_1, ack => convTranspose_CP_814_elements(88)); -- 
    -- CP-element group 89:  transition  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	86 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (6) 
      -- CP-element group 89: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_549_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_549_Sample/ra
      -- CP-element group 89: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_549_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_549_update_start_
      -- CP-element group 89: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_549_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_549_sample_completed_
      -- 
    ra_1525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_549_inst_ack_0, ack => convTranspose_CP_814_elements(89)); -- 
    cr_1529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(89), ack => RPIPE_ConvTranspose_input_pipe_549_inst_req_1); -- 
    -- CP-element group 90:  fork  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90: 	93 
    -- CP-element group 90:  members (9) 
      -- CP-element group 90: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_553_sample_start_
      -- CP-element group 90: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_549_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_553_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_549_Update/ca
      -- CP-element group 90: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_549_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_562_Sample/rr
      -- CP-element group 90: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_562_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_562_sample_start_
      -- CP-element group 90: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_553_Sample/rr
      -- 
    ca_1530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_549_inst_ack_1, ack => convTranspose_CP_814_elements(90)); -- 
    rr_1538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(90), ack => type_cast_553_inst_req_0); -- 
    rr_1552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(90), ack => RPIPE_ConvTranspose_input_pipe_562_inst_req_0); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_553_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_553_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_553_Sample/ra
      -- 
    ra_1539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_553_inst_ack_0, ack => convTranspose_CP_814_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	0 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	105 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_553_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_553_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_553_Update/$exit
      -- 
    ca_1544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_553_inst_ack_1, ack => convTranspose_CP_814_elements(92)); -- 
    -- CP-element group 93:  transition  input  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	90 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (6) 
      -- CP-element group 93: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_562_Update/$entry
      -- CP-element group 93: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_562_Update/cr
      -- CP-element group 93: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_562_Sample/ra
      -- CP-element group 93: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_562_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_562_update_start_
      -- CP-element group 93: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_562_sample_completed_
      -- 
    ra_1553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_562_inst_ack_0, ack => convTranspose_CP_814_elements(93)); -- 
    cr_1557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(93), ack => RPIPE_ConvTranspose_input_pipe_562_inst_req_1); -- 
    -- CP-element group 94:  fork  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94: 	97 
    -- CP-element group 94:  members (9) 
      -- CP-element group 94: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_574_Sample/rr
      -- CP-element group 94: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_574_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_566_Sample/rr
      -- CP-element group 94: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_566_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_574_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_566_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_562_Update/ca
      -- CP-element group 94: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_562_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_562_update_completed_
      -- 
    ca_1558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_562_inst_ack_1, ack => convTranspose_CP_814_elements(94)); -- 
    rr_1580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(94), ack => RPIPE_ConvTranspose_input_pipe_574_inst_req_0); -- 
    rr_1566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(94), ack => type_cast_566_inst_req_0); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_566_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_566_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_566_sample_completed_
      -- 
    ra_1567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_566_inst_ack_0, ack => convTranspose_CP_814_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	0 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	105 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_566_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_566_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_566_Update/$exit
      -- 
    ca_1572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_566_inst_ack_1, ack => convTranspose_CP_814_elements(96)); -- 
    -- CP-element group 97:  transition  input  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	94 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (6) 
      -- CP-element group 97: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_574_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_574_Update/$entry
      -- CP-element group 97: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_574_Sample/ra
      -- CP-element group 97: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_574_update_start_
      -- CP-element group 97: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_574_Update/cr
      -- CP-element group 97: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_574_Sample/$exit
      -- 
    ra_1581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_574_inst_ack_0, ack => convTranspose_CP_814_elements(97)); -- 
    cr_1585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(97), ack => RPIPE_ConvTranspose_input_pipe_574_inst_req_1); -- 
    -- CP-element group 98:  fork  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98: 	101 
    -- CP-element group 98:  members (9) 
      -- CP-element group 98: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_578_Sample/rr
      -- CP-element group 98: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_587_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_587_Sample/rr
      -- CP-element group 98: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_574_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_574_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_574_Update/ca
      -- CP-element group 98: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_578_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_587_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_578_sample_start_
      -- 
    ca_1586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_574_inst_ack_1, ack => convTranspose_CP_814_elements(98)); -- 
    rr_1594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(98), ack => type_cast_578_inst_req_0); -- 
    rr_1608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(98), ack => RPIPE_ConvTranspose_input_pipe_587_inst_req_0); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_578_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_578_Sample/ra
      -- CP-element group 99: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_578_sample_completed_
      -- 
    ra_1595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_578_inst_ack_0, ack => convTranspose_CP_814_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	0 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	105 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_578_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_578_Update/ca
      -- CP-element group 100: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_578_Update/$exit
      -- 
    ca_1600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_578_inst_ack_1, ack => convTranspose_CP_814_elements(100)); -- 
    -- CP-element group 101:  transition  input  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	98 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (6) 
      -- CP-element group 101: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_587_Sample/ra
      -- CP-element group 101: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_587_Update/$entry
      -- CP-element group 101: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_587_Update/cr
      -- CP-element group 101: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_587_update_start_
      -- CP-element group 101: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_587_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_587_sample_completed_
      -- 
    ra_1609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_587_inst_ack_0, ack => convTranspose_CP_814_elements(101)); -- 
    cr_1613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(101), ack => RPIPE_ConvTranspose_input_pipe_587_inst_req_1); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (6) 
      -- CP-element group 102: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_587_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_587_Update/ca
      -- CP-element group 102: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/RPIPE_ConvTranspose_input_pipe_587_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_591_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_591_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_591_Sample/$entry
      -- 
    ca_1614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_587_inst_ack_1, ack => convTranspose_CP_814_elements(102)); -- 
    rr_1622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(102), ack => type_cast_591_inst_req_0); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_591_Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_591_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_591_sample_completed_
      -- 
    ra_1623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_591_inst_ack_0, ack => convTranspose_CP_814_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	0 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_591_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_591_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/type_cast_591_update_completed_
      -- 
    ca_1628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_591_inst_ack_1, ack => convTranspose_CP_814_elements(104)); -- 
    -- CP-element group 105:  join  fork  transition  place  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	32 
    -- CP-element group 105: 	52 
    -- CP-element group 105: 	36 
    -- CP-element group 105: 	48 
    -- CP-element group 105: 	44 
    -- CP-element group 105: 	40 
    -- CP-element group 105: 	72 
    -- CP-element group 105: 	56 
    -- CP-element group 105: 	64 
    -- CP-element group 105: 	60 
    -- CP-element group 105: 	68 
    -- CP-element group 105: 	80 
    -- CP-element group 105: 	96 
    -- CP-element group 105: 	88 
    -- CP-element group 105: 	100 
    -- CP-element group 105: 	76 
    -- CP-element group 105: 	84 
    -- CP-element group 105: 	104 
    -- CP-element group 105: 	92 
    -- CP-element group 105: 	4 
    -- CP-element group 105: 	8 
    -- CP-element group 105: 	12 
    -- CP-element group 105: 	16 
    -- CP-element group 105: 	20 
    -- CP-element group 105: 	24 
    -- CP-element group 105: 	28 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	118 
    -- CP-element group 105: 	119 
    -- CP-element group 105: 	109 
    -- CP-element group 105: 	110 
    -- CP-element group 105: 	111 
    -- CP-element group 105: 	112 
    -- CP-element group 105: 	113 
    -- CP-element group 105: 	114 
    -- CP-element group 105: 	115 
    -- CP-element group 105: 	116 
    -- CP-element group 105: 	117 
    -- CP-element group 105: 	106 
    -- CP-element group 105: 	107 
    -- CP-element group 105: 	108 
    -- CP-element group 105:  members (46) 
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_609_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667__entry__
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597__exit__
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_641_Sample/rr
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_627_Sample/rr
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_641_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_605_Update/cr
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_605_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_627_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_641_Update/cr
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_623_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_623_Update/cr
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_274_to_assign_stmt_597/$exit
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_609_Sample/rr
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_609_Update/cr
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_609_update_start_
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_609_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_645_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_609_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_641_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_623_Sample/rr
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_623_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_645_update_start_
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_645_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_645_Sample/rr
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_627_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_645_Update/cr
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_627_Update/cr
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_641_update_start_
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_623_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_645_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_627_update_start_
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_623_update_start_
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_641_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_627_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_605_Sample/rr
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_605_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_605_update_start_
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_605_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_601_Update/cr
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_601_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_601_Sample/rr
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_601_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_601_update_start_
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_601_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/$entry
      -- 
    rr_1709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(105), ack => type_cast_641_inst_req_0); -- 
    rr_1695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(105), ack => type_cast_627_inst_req_0); -- 
    cr_1658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(105), ack => type_cast_605_inst_req_1); -- 
    cr_1714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(105), ack => type_cast_641_inst_req_1); -- 
    cr_1686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(105), ack => type_cast_623_inst_req_1); -- 
    rr_1667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(105), ack => type_cast_609_inst_req_0); -- 
    cr_1672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(105), ack => type_cast_609_inst_req_1); -- 
    rr_1681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(105), ack => type_cast_623_inst_req_0); -- 
    rr_1723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(105), ack => type_cast_645_inst_req_0); -- 
    cr_1728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(105), ack => type_cast_645_inst_req_1); -- 
    cr_1700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(105), ack => type_cast_627_inst_req_1); -- 
    rr_1653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(105), ack => type_cast_605_inst_req_0); -- 
    cr_1644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(105), ack => type_cast_601_inst_req_1); -- 
    rr_1639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(105), ack => type_cast_601_inst_req_0); -- 
    convTranspose_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 25) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1);
      constant place_markings: IntegerArray(0 to 25)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0);
      constant place_delays: IntegerArray(0 to 25) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 26); -- 
    begin -- 
      preds <= convTranspose_CP_814_elements(32) & convTranspose_CP_814_elements(52) & convTranspose_CP_814_elements(36) & convTranspose_CP_814_elements(48) & convTranspose_CP_814_elements(44) & convTranspose_CP_814_elements(40) & convTranspose_CP_814_elements(72) & convTranspose_CP_814_elements(56) & convTranspose_CP_814_elements(64) & convTranspose_CP_814_elements(60) & convTranspose_CP_814_elements(68) & convTranspose_CP_814_elements(80) & convTranspose_CP_814_elements(96) & convTranspose_CP_814_elements(88) & convTranspose_CP_814_elements(100) & convTranspose_CP_814_elements(76) & convTranspose_CP_814_elements(84) & convTranspose_CP_814_elements(104) & convTranspose_CP_814_elements(92) & convTranspose_CP_814_elements(4) & convTranspose_CP_814_elements(8) & convTranspose_CP_814_elements(12) & convTranspose_CP_814_elements(16) & convTranspose_CP_814_elements(20) & convTranspose_CP_814_elements(24) & convTranspose_CP_814_elements(28);
      gj_convTranspose_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 26, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_814_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_601_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_601_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_601_sample_completed_
      -- 
    ra_1640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_601_inst_ack_0, ack => convTranspose_CP_814_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	120 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_601_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_601_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_601_update_completed_
      -- 
    ca_1645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_601_inst_ack_1, ack => convTranspose_CP_814_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	105 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_605_Sample/ra
      -- CP-element group 108: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_605_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_605_sample_completed_
      -- 
    ra_1654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_605_inst_ack_0, ack => convTranspose_CP_814_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	105 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	120 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_605_Update/ca
      -- CP-element group 109: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_605_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_605_update_completed_
      -- 
    ca_1659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_605_inst_ack_1, ack => convTranspose_CP_814_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	105 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_609_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_609_Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_609_sample_completed_
      -- 
    ra_1668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_609_inst_ack_0, ack => convTranspose_CP_814_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	105 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	120 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_609_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_609_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_609_update_completed_
      -- 
    ca_1673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_609_inst_ack_1, ack => convTranspose_CP_814_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	105 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_623_Sample/ra
      -- CP-element group 112: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_623_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_623_sample_completed_
      -- 
    ra_1682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_623_inst_ack_0, ack => convTranspose_CP_814_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	105 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	120 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_623_Update/ca
      -- CP-element group 113: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_623_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_623_update_completed_
      -- 
    ca_1687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_623_inst_ack_1, ack => convTranspose_CP_814_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	105 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_627_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_627_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_627_sample_completed_
      -- 
    ra_1696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_627_inst_ack_0, ack => convTranspose_CP_814_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	105 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	120 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_627_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_627_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_627_Update/ca
      -- 
    ca_1701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_627_inst_ack_1, ack => convTranspose_CP_814_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	105 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_641_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_641_Sample/ra
      -- CP-element group 116: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_641_sample_completed_
      -- 
    ra_1710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_641_inst_ack_0, ack => convTranspose_CP_814_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	105 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	120 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_641_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_641_Update/ca
      -- CP-element group 117: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_641_update_completed_
      -- 
    ca_1715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_641_inst_ack_1, ack => convTranspose_CP_814_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	105 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_645_sample_completed_
      -- CP-element group 118: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_645_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_645_Sample/ra
      -- 
    ra_1724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_645_inst_ack_0, ack => convTranspose_CP_814_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	105 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_645_Update/ca
      -- CP-element group 119: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_645_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/type_cast_645_Update/$exit
      -- 
    ca_1729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_645_inst_ack_1, ack => convTranspose_CP_814_elements(119)); -- 
    -- CP-element group 120:  branch  join  transition  place  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: 	109 
    -- CP-element group 120: 	111 
    -- CP-element group 120: 	113 
    -- CP-element group 120: 	115 
    -- CP-element group 120: 	117 
    -- CP-element group 120: 	107 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (10) 
      -- CP-element group 120: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667__exit__
      -- CP-element group 120: 	 branch_block_stmt_271/if_stmt_668_eval_test/$entry
      -- CP-element group 120: 	 branch_block_stmt_271/if_stmt_668_eval_test/$exit
      -- CP-element group 120: 	 branch_block_stmt_271/if_stmt_668_eval_test/branch_req
      -- CP-element group 120: 	 branch_block_stmt_271/if_stmt_668_dead_link/$entry
      -- CP-element group 120: 	 branch_block_stmt_271/if_stmt_668__entry__
      -- CP-element group 120: 	 branch_block_stmt_271/R_cmp376_669_place
      -- CP-element group 120: 	 branch_block_stmt_271/if_stmt_668_else_link/$entry
      -- CP-element group 120: 	 branch_block_stmt_271/assign_stmt_602_to_assign_stmt_667/$exit
      -- CP-element group 120: 	 branch_block_stmt_271/if_stmt_668_if_link/$entry
      -- 
    branch_req_1737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(120), ack => if_stmt_668_branch_req_0); -- 
    convTranspose_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convTranspose_CP_814_elements(119) & convTranspose_CP_814_elements(109) & convTranspose_CP_814_elements(111) & convTranspose_CP_814_elements(113) & convTranspose_CP_814_elements(115) & convTranspose_CP_814_elements(117) & convTranspose_CP_814_elements(107);
      gj_convTranspose_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_814_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121: 	124 
    -- CP-element group 121:  members (18) 
      -- CP-element group 121: 	 branch_block_stmt_271/assign_stmt_680_to_assign_stmt_709/type_cast_695_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_271/assign_stmt_680_to_assign_stmt_709/type_cast_695_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_271/assign_stmt_680_to_assign_stmt_709/type_cast_695_update_start_
      -- CP-element group 121: 	 branch_block_stmt_271/assign_stmt_680_to_assign_stmt_709/type_cast_695_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_271/assign_stmt_680_to_assign_stmt_709/type_cast_695_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_271/assign_stmt_680_to_assign_stmt_709/type_cast_695_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_271/assign_stmt_680_to_assign_stmt_709__entry__
      -- CP-element group 121: 	 branch_block_stmt_271/merge_stmt_674__exit__
      -- CP-element group 121: 	 branch_block_stmt_271/entry_bbx_xnph378
      -- CP-element group 121: 	 branch_block_stmt_271/if_stmt_668_if_link/if_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_271/if_stmt_668_if_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_271/assign_stmt_680_to_assign_stmt_709/$entry
      -- CP-element group 121: 	 branch_block_stmt_271/merge_stmt_674_PhiAck/dummy
      -- CP-element group 121: 	 branch_block_stmt_271/merge_stmt_674_PhiAck/$exit
      -- CP-element group 121: 	 branch_block_stmt_271/merge_stmt_674_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_271/entry_bbx_xnph378_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_271/entry_bbx_xnph378_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_271/merge_stmt_674_PhiReqMerge
      -- 
    if_choice_transition_1742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_668_branch_ack_1, ack => convTranspose_CP_814_elements(121)); -- 
    cr_1764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(121), ack => type_cast_695_inst_req_1); -- 
    rr_1759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(121), ack => type_cast_695_inst_req_0); -- 
    -- CP-element group 122:  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	230 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_271/entry_forx_xend
      -- CP-element group 122: 	 branch_block_stmt_271/if_stmt_668_else_link/else_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_271/if_stmt_668_else_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_271/entry_forx_xend_PhiReq/$exit
      -- CP-element group 122: 	 branch_block_stmt_271/entry_forx_xend_PhiReq/$entry
      -- 
    else_choice_transition_1746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_668_branch_ack_0, ack => convTranspose_CP_814_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_271/assign_stmt_680_to_assign_stmt_709/type_cast_695_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_271/assign_stmt_680_to_assign_stmt_709/type_cast_695_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_271/assign_stmt_680_to_assign_stmt_709/type_cast_695_Sample/ra
      -- 
    ra_1760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_695_inst_ack_0, ack => convTranspose_CP_814_elements(123)); -- 
    -- CP-element group 124:  transition  place  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	121 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	224 
    -- CP-element group 124:  members (9) 
      -- CP-element group 124: 	 branch_block_stmt_271/assign_stmt_680_to_assign_stmt_709/type_cast_695_Update/ca
      -- CP-element group 124: 	 branch_block_stmt_271/assign_stmt_680_to_assign_stmt_709/type_cast_695_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_271/assign_stmt_680_to_assign_stmt_709/type_cast_695_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_271/bbx_xnph378_forx_xbody_PhiReq/phi_stmt_712/$entry
      -- CP-element group 124: 	 branch_block_stmt_271/bbx_xnph378_forx_xbody_PhiReq/$entry
      -- CP-element group 124: 	 branch_block_stmt_271/bbx_xnph378_forx_xbody
      -- CP-element group 124: 	 branch_block_stmt_271/assign_stmt_680_to_assign_stmt_709__exit__
      -- CP-element group 124: 	 branch_block_stmt_271/assign_stmt_680_to_assign_stmt_709/$exit
      -- CP-element group 124: 	 branch_block_stmt_271/bbx_xnph378_forx_xbody_PhiReq/phi_stmt_712/phi_stmt_712_sources/$entry
      -- 
    ca_1765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_695_inst_ack_1, ack => convTranspose_CP_814_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	229 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	164 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_final_index_sum_regn_sample_complete
      -- CP-element group 125: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_final_index_sum_regn_Sample/ack
      -- CP-element group 125: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_final_index_sum_regn_Sample/$exit
      -- 
    ack_1794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_724_index_offset_ack_0, ack => convTranspose_CP_814_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	229 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (11) 
      -- CP-element group 126: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_base_plus_offset/$entry
      -- CP-element group 126: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_final_index_sum_regn_Update/ack
      -- CP-element group 126: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/addr_of_725_request/$entry
      -- CP-element group 126: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_base_plus_offset/$exit
      -- CP-element group 126: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/addr_of_725_request/req
      -- CP-element group 126: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/addr_of_725_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_base_plus_offset/sum_rename_req
      -- CP-element group 126: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_base_plus_offset/sum_rename_ack
      -- CP-element group 126: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_final_index_sum_regn_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_offset_calculated
      -- CP-element group 126: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_root_address_calculated
      -- 
    ack_1799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_724_index_offset_ack_1, ack => convTranspose_CP_814_elements(126)); -- 
    req_1808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(126), ack => addr_of_725_final_reg_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/addr_of_725_request/ack
      -- CP-element group 127: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/addr_of_725_request/$exit
      -- CP-element group 127: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/addr_of_725_sample_completed_
      -- 
    ack_1809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_725_final_reg_ack_0, ack => convTranspose_CP_814_elements(127)); -- 
    -- CP-element group 128:  fork  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	229 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	161 
    -- CP-element group 128:  members (19) 
      -- CP-element group 128: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/addr_of_725_complete/$exit
      -- CP-element group 128: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/addr_of_725_complete/ack
      -- CP-element group 128: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/addr_of_725_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_base_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_word_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_root_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_base_address_resized
      -- CP-element group 128: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_base_addr_resize/$entry
      -- CP-element group 128: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_base_addr_resize/$exit
      -- CP-element group 128: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_base_addr_resize/base_resize_req
      -- CP-element group 128: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_base_addr_resize/base_resize_ack
      -- CP-element group 128: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_base_plus_offset/$entry
      -- CP-element group 128: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_base_plus_offset/$exit
      -- CP-element group 128: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_base_plus_offset/sum_rename_req
      -- CP-element group 128: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_base_plus_offset/sum_rename_ack
      -- CP-element group 128: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_word_addrgen/$entry
      -- CP-element group 128: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_word_addrgen/$exit
      -- CP-element group 128: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_word_addrgen/root_register_req
      -- CP-element group 128: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_word_addrgen/root_register_ack
      -- 
    ack_1814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_725_final_reg_ack_1, ack => convTranspose_CP_814_elements(128)); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	229 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_728_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_728_Sample/ra
      -- CP-element group 129: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_728_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_728_Update/cr
      -- CP-element group 129: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_728_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_728_update_start_
      -- 
    ra_1823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_728_inst_ack_0, ack => convTranspose_CP_814_elements(129)); -- 
    cr_1827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(129), ack => RPIPE_ConvTranspose_input_pipe_728_inst_req_1); -- 
    -- CP-element group 130:  fork  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (9) 
      -- CP-element group 130: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_728_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_728_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_741_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_741_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_728_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_732_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_732_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_741_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_732_Sample/rr
      -- 
    ca_1828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_728_inst_ack_1, ack => convTranspose_CP_814_elements(130)); -- 
    rr_1836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(130), ack => type_cast_732_inst_req_0); -- 
    rr_1850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(130), ack => RPIPE_ConvTranspose_input_pipe_741_inst_req_0); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_732_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_732_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_732_Sample/ra
      -- 
    ra_1837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_732_inst_ack_0, ack => convTranspose_CP_814_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	229 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	161 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_732_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_732_Update/ca
      -- CP-element group 132: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_732_Update/$exit
      -- 
    ca_1842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_732_inst_ack_1, ack => convTranspose_CP_814_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_741_update_start_
      -- CP-element group 133: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_741_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_741_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_741_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_741_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_741_Update/cr
      -- 
    ra_1851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_741_inst_ack_0, ack => convTranspose_CP_814_elements(133)); -- 
    cr_1855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(133), ack => RPIPE_ConvTranspose_input_pipe_741_inst_req_1); -- 
    -- CP-element group 134:  fork  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (9) 
      -- CP-element group 134: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_741_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_745_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_741_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_745_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_741_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_759_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_759_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_745_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_759_Sample/rr
      -- 
    ca_1856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_741_inst_ack_1, ack => convTranspose_CP_814_elements(134)); -- 
    rr_1864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(134), ack => type_cast_745_inst_req_0); -- 
    rr_1878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(134), ack => RPIPE_ConvTranspose_input_pipe_759_inst_req_0); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_745_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_745_Sample/ra
      -- CP-element group 135: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_745_Sample/$exit
      -- 
    ra_1865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_745_inst_ack_0, ack => convTranspose_CP_814_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	229 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	161 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_745_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_745_Update/ca
      -- CP-element group 136: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_745_update_completed_
      -- 
    ca_1870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_745_inst_ack_1, ack => convTranspose_CP_814_elements(136)); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_759_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_759_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_759_update_start_
      -- CP-element group 137: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_759_Sample/ra
      -- CP-element group 137: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_759_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_759_Update/cr
      -- 
    ra_1879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_759_inst_ack_0, ack => convTranspose_CP_814_elements(137)); -- 
    cr_1883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(137), ack => RPIPE_ConvTranspose_input_pipe_759_inst_req_1); -- 
    -- CP-element group 138:  fork  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138: 	141 
    -- CP-element group 138:  members (9) 
      -- CP-element group 138: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_759_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_759_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_759_Update/ca
      -- CP-element group 138: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_763_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_763_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_763_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_777_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_777_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_777_Sample/rr
      -- 
    ca_1884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_759_inst_ack_1, ack => convTranspose_CP_814_elements(138)); -- 
    rr_1892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(138), ack => type_cast_763_inst_req_0); -- 
    rr_1906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(138), ack => RPIPE_ConvTranspose_input_pipe_777_inst_req_0); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_763_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_763_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_763_Sample/ra
      -- 
    ra_1893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_763_inst_ack_0, ack => convTranspose_CP_814_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	229 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	161 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_763_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_763_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_763_Update/ca
      -- 
    ca_1898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_763_inst_ack_1, ack => convTranspose_CP_814_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	138 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (6) 
      -- CP-element group 141: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_777_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_777_update_start_
      -- CP-element group 141: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_777_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_777_Sample/ra
      -- CP-element group 141: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_777_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_777_Update/cr
      -- 
    ra_1907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_777_inst_ack_0, ack => convTranspose_CP_814_elements(141)); -- 
    cr_1911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(141), ack => RPIPE_ConvTranspose_input_pipe_777_inst_req_1); -- 
    -- CP-element group 142:  fork  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	145 
    -- CP-element group 142:  members (9) 
      -- CP-element group 142: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_777_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_777_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_777_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_781_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_781_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_781_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_795_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_795_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_795_Sample/rr
      -- 
    ca_1912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_777_inst_ack_1, ack => convTranspose_CP_814_elements(142)); -- 
    rr_1920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(142), ack => type_cast_781_inst_req_0); -- 
    rr_1934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(142), ack => RPIPE_ConvTranspose_input_pipe_795_inst_req_0); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_781_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_781_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_781_Sample/ra
      -- 
    ra_1921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_781_inst_ack_0, ack => convTranspose_CP_814_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	229 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	161 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_781_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_781_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_781_Update/ca
      -- 
    ca_1926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_781_inst_ack_1, ack => convTranspose_CP_814_elements(144)); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	142 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_795_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_795_update_start_
      -- CP-element group 145: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_795_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_795_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_795_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_795_Update/cr
      -- 
    ra_1935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_795_inst_ack_0, ack => convTranspose_CP_814_elements(145)); -- 
    cr_1939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(145), ack => RPIPE_ConvTranspose_input_pipe_795_inst_req_1); -- 
    -- CP-element group 146:  fork  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	149 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_795_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_795_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_795_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_799_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_799_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_799_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_813_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_813_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_813_Sample/rr
      -- 
    ca_1940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_795_inst_ack_1, ack => convTranspose_CP_814_elements(146)); -- 
    rr_1962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(146), ack => RPIPE_ConvTranspose_input_pipe_813_inst_req_0); -- 
    rr_1948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(146), ack => type_cast_799_inst_req_0); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_799_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_799_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_799_Sample/ra
      -- 
    ra_1949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_799_inst_ack_0, ack => convTranspose_CP_814_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	229 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	161 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_799_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_799_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_799_Update/ca
      -- 
    ca_1954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_799_inst_ack_1, ack => convTranspose_CP_814_elements(148)); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	146 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_813_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_813_update_start_
      -- CP-element group 149: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_813_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_813_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_813_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_813_Update/cr
      -- 
    ra_1963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_813_inst_ack_0, ack => convTranspose_CP_814_elements(149)); -- 
    cr_1967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(149), ack => RPIPE_ConvTranspose_input_pipe_813_inst_req_1); -- 
    -- CP-element group 150:  fork  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (9) 
      -- CP-element group 150: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_813_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_813_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_813_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_817_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_817_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_817_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_831_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_831_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_831_Sample/rr
      -- 
    ca_1968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_813_inst_ack_1, ack => convTranspose_CP_814_elements(150)); -- 
    rr_1976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(150), ack => type_cast_817_inst_req_0); -- 
    rr_1990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(150), ack => RPIPE_ConvTranspose_input_pipe_831_inst_req_0); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_817_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_817_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_817_Sample/ra
      -- 
    ra_1977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_817_inst_ack_0, ack => convTranspose_CP_814_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	229 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	161 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_817_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_817_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_817_Update/ca
      -- 
    ca_1982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_817_inst_ack_1, ack => convTranspose_CP_814_elements(152)); -- 
    -- CP-element group 153:  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	150 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (6) 
      -- CP-element group 153: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_831_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_831_update_start_
      -- CP-element group 153: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_831_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_831_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_831_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_831_Update/cr
      -- 
    ra_1991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_831_inst_ack_0, ack => convTranspose_CP_814_elements(153)); -- 
    cr_1995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(153), ack => RPIPE_ConvTranspose_input_pipe_831_inst_req_1); -- 
    -- CP-element group 154:  fork  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154: 	157 
    -- CP-element group 154:  members (9) 
      -- CP-element group 154: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_831_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_831_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_831_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_835_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_835_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_835_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_849_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_849_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_849_Sample/rr
      -- 
    ca_1996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_831_inst_ack_1, ack => convTranspose_CP_814_elements(154)); -- 
    rr_2004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(154), ack => type_cast_835_inst_req_0); -- 
    rr_2018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(154), ack => RPIPE_ConvTranspose_input_pipe_849_inst_req_0); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_835_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_835_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_835_Sample/ra
      -- 
    ra_2005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_835_inst_ack_0, ack => convTranspose_CP_814_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	229 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	161 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_835_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_835_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_835_Update/ca
      -- 
    ca_2010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_835_inst_ack_1, ack => convTranspose_CP_814_elements(156)); -- 
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_849_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_849_update_start_
      -- CP-element group 157: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_849_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_849_Sample/ra
      -- CP-element group 157: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_849_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_849_Update/cr
      -- 
    ra_2019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_849_inst_ack_0, ack => convTranspose_CP_814_elements(157)); -- 
    cr_2023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(157), ack => RPIPE_ConvTranspose_input_pipe_849_inst_req_1); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_849_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_849_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_849_Update/ca
      -- CP-element group 158: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_853_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_853_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_853_Sample/rr
      -- 
    ca_2024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_849_inst_ack_1, ack => convTranspose_CP_814_elements(158)); -- 
    rr_2032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(158), ack => type_cast_853_inst_req_0); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_853_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_853_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_853_Sample/ra
      -- 
    ra_2033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_853_inst_ack_0, ack => convTranspose_CP_814_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	229 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_853_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_853_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_853_Update/ca
      -- 
    ca_2038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_853_inst_ack_1, ack => convTranspose_CP_814_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	148 
    -- CP-element group 161: 	152 
    -- CP-element group 161: 	156 
    -- CP-element group 161: 	160 
    -- CP-element group 161: 	132 
    -- CP-element group 161: 	128 
    -- CP-element group 161: 	144 
    -- CP-element group 161: 	140 
    -- CP-element group 161: 	136 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (9) 
      -- CP-element group 161: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_Sample/ptr_deref_861_Split/$entry
      -- CP-element group 161: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_Sample/ptr_deref_861_Split/$exit
      -- CP-element group 161: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_Sample/ptr_deref_861_Split/split_req
      -- CP-element group 161: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_Sample/ptr_deref_861_Split/split_ack
      -- CP-element group 161: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_Sample/word_access_start/$entry
      -- CP-element group 161: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_Sample/word_access_start/word_0/$entry
      -- CP-element group 161: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_Sample/word_access_start/word_0/rr
      -- 
    rr_2076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(161), ack => ptr_deref_861_store_0_req_0); -- 
    convTranspose_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_814_elements(148) & convTranspose_CP_814_elements(152) & convTranspose_CP_814_elements(156) & convTranspose_CP_814_elements(160) & convTranspose_CP_814_elements(132) & convTranspose_CP_814_elements(128) & convTranspose_CP_814_elements(144) & convTranspose_CP_814_elements(140) & convTranspose_CP_814_elements(136);
      gj_convTranspose_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_814_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_Sample/word_access_start/$exit
      -- CP-element group 162: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_Sample/word_access_start/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_Sample/word_access_start/word_0/ra
      -- 
    ra_2077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_861_store_0_ack_0, ack => convTranspose_CP_814_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	229 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_Update/word_access_complete/$exit
      -- CP-element group 163: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_Update/word_access_complete/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_Update/word_access_complete/word_0/ca
      -- 
    ca_2088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_861_store_0_ack_1, ack => convTranspose_CP_814_elements(163)); -- 
    -- CP-element group 164:  branch  join  transition  place  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: 	125 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (10) 
      -- CP-element group 164: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/$exit
      -- CP-element group 164: 	 branch_block_stmt_271/if_stmt_875__entry__
      -- CP-element group 164: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874__exit__
      -- CP-element group 164: 	 branch_block_stmt_271/if_stmt_875_dead_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_271/if_stmt_875_eval_test/$entry
      -- CP-element group 164: 	 branch_block_stmt_271/if_stmt_875_eval_test/$exit
      -- CP-element group 164: 	 branch_block_stmt_271/if_stmt_875_eval_test/branch_req
      -- CP-element group 164: 	 branch_block_stmt_271/R_exitcond2_876_place
      -- CP-element group 164: 	 branch_block_stmt_271/if_stmt_875_if_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_271/if_stmt_875_else_link/$entry
      -- 
    branch_req_2096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(164), ack => if_stmt_875_branch_req_0); -- 
    convTranspose_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_814_elements(163) & convTranspose_CP_814_elements(125);
      gj_convTranspose_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_814_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  merge  transition  place  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	230 
    -- CP-element group 165:  members (13) 
      -- CP-element group 165: 	 branch_block_stmt_271/forx_xendx_xloopexit_forx_xend
      -- CP-element group 165: 	 branch_block_stmt_271/merge_stmt_881__exit__
      -- CP-element group 165: 	 branch_block_stmt_271/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_271/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_271/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_271/if_stmt_875_if_link/$exit
      -- CP-element group 165: 	 branch_block_stmt_271/if_stmt_875_if_link/if_choice_transition
      -- CP-element group 165: 	 branch_block_stmt_271/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 165: 	 branch_block_stmt_271/merge_stmt_881_PhiAck/dummy
      -- CP-element group 165: 	 branch_block_stmt_271/merge_stmt_881_PhiAck/$exit
      -- CP-element group 165: 	 branch_block_stmt_271/merge_stmt_881_PhiAck/$entry
      -- CP-element group 165: 	 branch_block_stmt_271/merge_stmt_881_PhiReqMerge
      -- CP-element group 165: 	 branch_block_stmt_271/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- 
    if_choice_transition_2101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_875_branch_ack_1, ack => convTranspose_CP_814_elements(165)); -- 
    -- CP-element group 166:  fork  transition  place  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	225 
    -- CP-element group 166: 	226 
    -- CP-element group 166:  members (12) 
      -- CP-element group 166: 	 branch_block_stmt_271/forx_xbody_forx_xbody_PhiReq/phi_stmt_712/phi_stmt_712_sources/type_cast_718/SplitProtocol/Update/cr
      -- CP-element group 166: 	 branch_block_stmt_271/forx_xbody_forx_xbody_PhiReq/phi_stmt_712/phi_stmt_712_sources/type_cast_718/SplitProtocol/Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_271/forx_xbody_forx_xbody_PhiReq/phi_stmt_712/phi_stmt_712_sources/type_cast_718/SplitProtocol/Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_271/forx_xbody_forx_xbody_PhiReq/phi_stmt_712/phi_stmt_712_sources/type_cast_718/SplitProtocol/Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_271/forx_xbody_forx_xbody_PhiReq/phi_stmt_712/phi_stmt_712_sources/type_cast_718/SplitProtocol/$entry
      -- CP-element group 166: 	 branch_block_stmt_271/forx_xbody_forx_xbody_PhiReq/phi_stmt_712/phi_stmt_712_sources/type_cast_718/$entry
      -- CP-element group 166: 	 branch_block_stmt_271/forx_xbody_forx_xbody_PhiReq/phi_stmt_712/phi_stmt_712_sources/$entry
      -- CP-element group 166: 	 branch_block_stmt_271/if_stmt_875_else_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_271/if_stmt_875_else_link/else_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_271/forx_xbody_forx_xbody
      -- CP-element group 166: 	 branch_block_stmt_271/forx_xbody_forx_xbody_PhiReq/phi_stmt_712/$entry
      -- CP-element group 166: 	 branch_block_stmt_271/forx_xbody_forx_xbody_PhiReq/$entry
      -- 
    else_choice_transition_2105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_875_branch_ack_0, ack => convTranspose_CP_814_elements(166)); -- 
    cr_2755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(166), ack => type_cast_718_inst_req_1); -- 
    rr_2750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(166), ack => type_cast_718_inst_req_0); -- 
    -- CP-element group 167:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	230 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167: 	170 
    -- CP-element group 167:  members (18) 
      -- CP-element group 167: 	 branch_block_stmt_271/assign_stmt_902_to_assign_stmt_947__entry__
      -- CP-element group 167: 	 branch_block_stmt_271/merge_stmt_897__exit__
      -- CP-element group 167: 	 branch_block_stmt_271/forx_xend_bbx_xnph374_PhiReq/$exit
      -- CP-element group 167: 	 branch_block_stmt_271/forx_xend_bbx_xnph374_PhiReq/$entry
      -- CP-element group 167: 	 branch_block_stmt_271/merge_stmt_897_PhiAck/dummy
      -- CP-element group 167: 	 branch_block_stmt_271/merge_stmt_897_PhiAck/$exit
      -- CP-element group 167: 	 branch_block_stmt_271/if_stmt_891_if_link/$exit
      -- CP-element group 167: 	 branch_block_stmt_271/if_stmt_891_if_link/if_choice_transition
      -- CP-element group 167: 	 branch_block_stmt_271/forx_xend_bbx_xnph374
      -- CP-element group 167: 	 branch_block_stmt_271/assign_stmt_902_to_assign_stmt_947/$entry
      -- CP-element group 167: 	 branch_block_stmt_271/assign_stmt_902_to_assign_stmt_947/type_cast_933_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_271/assign_stmt_902_to_assign_stmt_947/type_cast_933_update_start_
      -- CP-element group 167: 	 branch_block_stmt_271/assign_stmt_902_to_assign_stmt_947/type_cast_933_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_271/assign_stmt_902_to_assign_stmt_947/type_cast_933_Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_271/assign_stmt_902_to_assign_stmt_947/type_cast_933_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_271/assign_stmt_902_to_assign_stmt_947/type_cast_933_Update/cr
      -- CP-element group 167: 	 branch_block_stmt_271/merge_stmt_897_PhiAck/$entry
      -- CP-element group 167: 	 branch_block_stmt_271/merge_stmt_897_PhiReqMerge
      -- 
    if_choice_transition_2123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_891_branch_ack_1, ack => convTranspose_CP_814_elements(167)); -- 
    rr_2140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(167), ack => type_cast_933_inst_req_0); -- 
    cr_2145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(167), ack => type_cast_933_inst_req_1); -- 
    -- CP-element group 168:  transition  place  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	230 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	237 
    -- CP-element group 168:  members (5) 
      -- CP-element group 168: 	 branch_block_stmt_271/if_stmt_891_else_link/$exit
      -- CP-element group 168: 	 branch_block_stmt_271/if_stmt_891_else_link/else_choice_transition
      -- CP-element group 168: 	 branch_block_stmt_271/forx_xend_forx_xend220
      -- CP-element group 168: 	 branch_block_stmt_271/forx_xend_forx_xend220_PhiReq/$entry
      -- CP-element group 168: 	 branch_block_stmt_271/forx_xend_forx_xend220_PhiReq/$exit
      -- 
    else_choice_transition_2127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_891_branch_ack_0, ack => convTranspose_CP_814_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_271/assign_stmt_902_to_assign_stmt_947/type_cast_933_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_271/assign_stmt_902_to_assign_stmt_947/type_cast_933_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_271/assign_stmt_902_to_assign_stmt_947/type_cast_933_Sample/ra
      -- 
    ra_2141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_933_inst_ack_0, ack => convTranspose_CP_814_elements(169)); -- 
    -- CP-element group 170:  transition  place  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	167 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	231 
    -- CP-element group 170:  members (9) 
      -- CP-element group 170: 	 branch_block_stmt_271/bbx_xnph374_forx_xbody214
      -- CP-element group 170: 	 branch_block_stmt_271/assign_stmt_902_to_assign_stmt_947__exit__
      -- CP-element group 170: 	 branch_block_stmt_271/bbx_xnph374_forx_xbody214_PhiReq/phi_stmt_950/phi_stmt_950_sources/$entry
      -- CP-element group 170: 	 branch_block_stmt_271/bbx_xnph374_forx_xbody214_PhiReq/phi_stmt_950/$entry
      -- CP-element group 170: 	 branch_block_stmt_271/bbx_xnph374_forx_xbody214_PhiReq/$entry
      -- CP-element group 170: 	 branch_block_stmt_271/assign_stmt_902_to_assign_stmt_947/$exit
      -- CP-element group 170: 	 branch_block_stmt_271/assign_stmt_902_to_assign_stmt_947/type_cast_933_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_271/assign_stmt_902_to_assign_stmt_947/type_cast_933_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_271/assign_stmt_902_to_assign_stmt_947/type_cast_933_Update/ca
      -- 
    ca_2146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_933_inst_ack_1, ack => convTranspose_CP_814_elements(170)); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	236 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_271/call_stmt_959_to_assign_stmt_970/call_stmt_959_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_271/call_stmt_959_to_assign_stmt_970/call_stmt_959_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_271/call_stmt_959_to_assign_stmt_970/call_stmt_959_Sample/cra
      -- 
    cra_2158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_959_call_ack_0, ack => convTranspose_CP_814_elements(171)); -- 
    -- CP-element group 172:  branch  transition  place  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	236 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (13) 
      -- CP-element group 172: 	 branch_block_stmt_271/if_stmt_971__entry__
      -- CP-element group 172: 	 branch_block_stmt_271/call_stmt_959_to_assign_stmt_970__exit__
      -- CP-element group 172: 	 branch_block_stmt_271/call_stmt_959_to_assign_stmt_970/$exit
      -- CP-element group 172: 	 branch_block_stmt_271/call_stmt_959_to_assign_stmt_970/call_stmt_959_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_271/call_stmt_959_to_assign_stmt_970/call_stmt_959_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_271/call_stmt_959_to_assign_stmt_970/call_stmt_959_Update/cca
      -- CP-element group 172: 	 branch_block_stmt_271/if_stmt_971_dead_link/$entry
      -- CP-element group 172: 	 branch_block_stmt_271/if_stmt_971_eval_test/$entry
      -- CP-element group 172: 	 branch_block_stmt_271/if_stmt_971_eval_test/$exit
      -- CP-element group 172: 	 branch_block_stmt_271/if_stmt_971_eval_test/branch_req
      -- CP-element group 172: 	 branch_block_stmt_271/R_exitcond_972_place
      -- CP-element group 172: 	 branch_block_stmt_271/if_stmt_971_if_link/$entry
      -- CP-element group 172: 	 branch_block_stmt_271/if_stmt_971_else_link/$entry
      -- 
    cca_2163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_959_call_ack_1, ack => convTranspose_CP_814_elements(172)); -- 
    branch_req_2171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(172), ack => if_stmt_971_branch_req_0); -- 
    -- CP-element group 173:  merge  transition  place  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	237 
    -- CP-element group 173:  members (13) 
      -- CP-element group 173: 	 branch_block_stmt_271/forx_xend220x_xloopexit_forx_xend220
      -- CP-element group 173: 	 branch_block_stmt_271/merge_stmt_977__exit__
      -- CP-element group 173: 	 branch_block_stmt_271/merge_stmt_977_PhiReqMerge
      -- CP-element group 173: 	 branch_block_stmt_271/merge_stmt_977_PhiAck/dummy
      -- CP-element group 173: 	 branch_block_stmt_271/forx_xbody214_forx_xend220x_xloopexit_PhiReq/$exit
      -- CP-element group 173: 	 branch_block_stmt_271/merge_stmt_977_PhiAck/$exit
      -- CP-element group 173: 	 branch_block_stmt_271/merge_stmt_977_PhiAck/$entry
      -- CP-element group 173: 	 branch_block_stmt_271/forx_xbody214_forx_xend220x_xloopexit_PhiReq/$entry
      -- CP-element group 173: 	 branch_block_stmt_271/if_stmt_971_if_link/$exit
      -- CP-element group 173: 	 branch_block_stmt_271/if_stmt_971_if_link/if_choice_transition
      -- CP-element group 173: 	 branch_block_stmt_271/forx_xbody214_forx_xend220x_xloopexit
      -- CP-element group 173: 	 branch_block_stmt_271/forx_xend220x_xloopexit_forx_xend220_PhiReq/$entry
      -- CP-element group 173: 	 branch_block_stmt_271/forx_xend220x_xloopexit_forx_xend220_PhiReq/$exit
      -- 
    if_choice_transition_2176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_971_branch_ack_1, ack => convTranspose_CP_814_elements(173)); -- 
    -- CP-element group 174:  fork  transition  place  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	232 
    -- CP-element group 174: 	233 
    -- CP-element group 174:  members (12) 
      -- CP-element group 174: 	 branch_block_stmt_271/forx_xbody214_forx_xbody214_PhiReq/phi_stmt_950/phi_stmt_950_sources/type_cast_956/SplitProtocol/Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_271/forx_xbody214_forx_xbody214_PhiReq/phi_stmt_950/phi_stmt_950_sources/type_cast_956/SplitProtocol/Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_271/forx_xbody214_forx_xbody214_PhiReq/phi_stmt_950/phi_stmt_950_sources/type_cast_956/SplitProtocol/Update/cr
      -- CP-element group 174: 	 branch_block_stmt_271/forx_xbody214_forx_xbody214_PhiReq/phi_stmt_950/phi_stmt_950_sources/type_cast_956/SplitProtocol/$entry
      -- CP-element group 174: 	 branch_block_stmt_271/forx_xbody214_forx_xbody214_PhiReq/phi_stmt_950/phi_stmt_950_sources/type_cast_956/$entry
      -- CP-element group 174: 	 branch_block_stmt_271/forx_xbody214_forx_xbody214_PhiReq/phi_stmt_950/phi_stmt_950_sources/type_cast_956/SplitProtocol/Update/$entry
      -- CP-element group 174: 	 branch_block_stmt_271/forx_xbody214_forx_xbody214_PhiReq/phi_stmt_950/phi_stmt_950_sources/$entry
      -- CP-element group 174: 	 branch_block_stmt_271/forx_xbody214_forx_xbody214_PhiReq/phi_stmt_950/$entry
      -- CP-element group 174: 	 branch_block_stmt_271/forx_xbody214_forx_xbody214_PhiReq/$entry
      -- CP-element group 174: 	 branch_block_stmt_271/if_stmt_971_else_link/$exit
      -- CP-element group 174: 	 branch_block_stmt_271/if_stmt_971_else_link/else_choice_transition
      -- CP-element group 174: 	 branch_block_stmt_271/forx_xbody214_forx_xbody214
      -- 
    else_choice_transition_2180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_971_branch_ack_0, ack => convTranspose_CP_814_elements(174)); -- 
    rr_2827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(174), ack => type_cast_956_inst_req_0); -- 
    cr_2832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(174), ack => type_cast_956_inst_req_1); -- 
    -- CP-element group 175:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	237 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175: 	178 
    -- CP-element group 175:  members (18) 
      -- CP-element group 175: 	 branch_block_stmt_271/merge_stmt_993__exit__
      -- CP-element group 175: 	 branch_block_stmt_271/assign_stmt_999_to_assign_stmt_1028__entry__
      -- CP-element group 175: 	 branch_block_stmt_271/if_stmt_987_if_link/$exit
      -- CP-element group 175: 	 branch_block_stmt_271/if_stmt_987_if_link/if_choice_transition
      -- CP-element group 175: 	 branch_block_stmt_271/forx_xend220_bbx_xnph
      -- CP-element group 175: 	 branch_block_stmt_271/assign_stmt_999_to_assign_stmt_1028/$entry
      -- CP-element group 175: 	 branch_block_stmt_271/assign_stmt_999_to_assign_stmt_1028/type_cast_1014_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_271/assign_stmt_999_to_assign_stmt_1028/type_cast_1014_update_start_
      -- CP-element group 175: 	 branch_block_stmt_271/assign_stmt_999_to_assign_stmt_1028/type_cast_1014_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_271/assign_stmt_999_to_assign_stmt_1028/type_cast_1014_Sample/rr
      -- CP-element group 175: 	 branch_block_stmt_271/assign_stmt_999_to_assign_stmt_1028/type_cast_1014_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_271/assign_stmt_999_to_assign_stmt_1028/type_cast_1014_Update/cr
      -- CP-element group 175: 	 branch_block_stmt_271/forx_xend220_bbx_xnph_PhiReq/$entry
      -- CP-element group 175: 	 branch_block_stmt_271/forx_xend220_bbx_xnph_PhiReq/$exit
      -- CP-element group 175: 	 branch_block_stmt_271/merge_stmt_993_PhiReqMerge
      -- CP-element group 175: 	 branch_block_stmt_271/merge_stmt_993_PhiAck/$entry
      -- CP-element group 175: 	 branch_block_stmt_271/merge_stmt_993_PhiAck/$exit
      -- CP-element group 175: 	 branch_block_stmt_271/merge_stmt_993_PhiAck/dummy
      -- 
    if_choice_transition_2198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_987_branch_ack_1, ack => convTranspose_CP_814_elements(175)); -- 
    rr_2215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(175), ack => type_cast_1014_inst_req_0); -- 
    cr_2220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(175), ack => type_cast_1014_inst_req_1); -- 
    -- CP-element group 176:  transition  place  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	237 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	244 
    -- CP-element group 176:  members (5) 
      -- CP-element group 176: 	 branch_block_stmt_271/if_stmt_987_else_link/$exit
      -- CP-element group 176: 	 branch_block_stmt_271/if_stmt_987_else_link/else_choice_transition
      -- CP-element group 176: 	 branch_block_stmt_271/forx_xend220_forx_xend235
      -- CP-element group 176: 	 branch_block_stmt_271/forx_xend220_forx_xend235_PhiReq/$entry
      -- CP-element group 176: 	 branch_block_stmt_271/forx_xend220_forx_xend235_PhiReq/$exit
      -- 
    else_choice_transition_2202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_987_branch_ack_0, ack => convTranspose_CP_814_elements(176)); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_271/assign_stmt_999_to_assign_stmt_1028/type_cast_1014_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_271/assign_stmt_999_to_assign_stmt_1028/type_cast_1014_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_271/assign_stmt_999_to_assign_stmt_1028/type_cast_1014_Sample/ra
      -- 
    ra_2216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1014_inst_ack_0, ack => convTranspose_CP_814_elements(177)); -- 
    -- CP-element group 178:  transition  place  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	175 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	238 
    -- CP-element group 178:  members (9) 
      -- CP-element group 178: 	 branch_block_stmt_271/bbx_xnph_forx_xbody228
      -- CP-element group 178: 	 branch_block_stmt_271/assign_stmt_999_to_assign_stmt_1028__exit__
      -- CP-element group 178: 	 branch_block_stmt_271/assign_stmt_999_to_assign_stmt_1028/$exit
      -- CP-element group 178: 	 branch_block_stmt_271/assign_stmt_999_to_assign_stmt_1028/type_cast_1014_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_271/assign_stmt_999_to_assign_stmt_1028/type_cast_1014_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_271/assign_stmt_999_to_assign_stmt_1028/type_cast_1014_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_271/bbx_xnph_forx_xbody228_PhiReq/$entry
      -- CP-element group 178: 	 branch_block_stmt_271/bbx_xnph_forx_xbody228_PhiReq/phi_stmt_1031/$entry
      -- CP-element group 178: 	 branch_block_stmt_271/bbx_xnph_forx_xbody228_PhiReq/phi_stmt_1031/phi_stmt_1031_sources/$entry
      -- 
    ca_2221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1014_inst_ack_1, ack => convTranspose_CP_814_elements(178)); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	243 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	185 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_final_index_sum_regn_sample_complete
      -- CP-element group 179: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_final_index_sum_regn_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_final_index_sum_regn_Sample/ack
      -- 
    ack_2250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1043_index_offset_ack_0, ack => convTranspose_CP_814_elements(179)); -- 
    -- CP-element group 180:  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	243 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (11) 
      -- CP-element group 180: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/addr_of_1044_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_root_address_calculated
      -- CP-element group 180: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_offset_calculated
      -- CP-element group 180: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_final_index_sum_regn_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_final_index_sum_regn_Update/ack
      -- CP-element group 180: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_base_plus_offset/$entry
      -- CP-element group 180: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_base_plus_offset/$exit
      -- CP-element group 180: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_base_plus_offset/sum_rename_req
      -- CP-element group 180: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_base_plus_offset/sum_rename_ack
      -- CP-element group 180: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/addr_of_1044_request/$entry
      -- CP-element group 180: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/addr_of_1044_request/req
      -- 
    ack_2255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1043_index_offset_ack_1, ack => convTranspose_CP_814_elements(180)); -- 
    req_2264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(180), ack => addr_of_1044_final_reg_req_0); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/addr_of_1044_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/addr_of_1044_request/$exit
      -- CP-element group 181: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/addr_of_1044_request/ack
      -- 
    ack_2265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1044_final_reg_ack_0, ack => convTranspose_CP_814_elements(181)); -- 
    -- CP-element group 182:  join  fork  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	243 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182:  members (28) 
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/addr_of_1044_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/addr_of_1044_complete/$exit
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/addr_of_1044_complete/ack
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_base_address_calculated
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_word_address_calculated
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_root_address_calculated
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_base_address_resized
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_base_addr_resize/$entry
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_base_addr_resize/$exit
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_base_addr_resize/base_resize_req
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_base_addr_resize/base_resize_ack
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_base_plus_offset/$entry
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_base_plus_offset/$exit
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_base_plus_offset/sum_rename_req
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_base_plus_offset/sum_rename_ack
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_word_addrgen/$entry
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_word_addrgen/$exit
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_word_addrgen/root_register_req
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_word_addrgen/root_register_ack
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_Sample/ptr_deref_1047_Split/$entry
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_Sample/ptr_deref_1047_Split/$exit
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_Sample/ptr_deref_1047_Split/split_req
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_Sample/ptr_deref_1047_Split/split_ack
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_Sample/word_access_start/$entry
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_Sample/word_access_start/word_0/$entry
      -- CP-element group 182: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_Sample/word_access_start/word_0/rr
      -- 
    ack_2270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1044_final_reg_ack_1, ack => convTranspose_CP_814_elements(182)); -- 
    rr_2308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(182), ack => ptr_deref_1047_store_0_req_0); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (5) 
      -- CP-element group 183: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_Sample/word_access_start/$exit
      -- CP-element group 183: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_Sample/word_access_start/word_0/$exit
      -- CP-element group 183: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_Sample/word_access_start/word_0/ra
      -- 
    ra_2309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1047_store_0_ack_0, ack => convTranspose_CP_814_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	243 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184:  members (5) 
      -- CP-element group 184: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_Update/word_access_complete/$exit
      -- CP-element group 184: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_Update/word_access_complete/word_0/$exit
      -- CP-element group 184: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_Update/word_access_complete/word_0/ca
      -- 
    ca_2320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1047_store_0_ack_1, ack => convTranspose_CP_814_elements(184)); -- 
    -- CP-element group 185:  branch  join  transition  place  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	179 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185: 	187 
    -- CP-element group 185:  members (10) 
      -- CP-element group 185: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061__exit__
      -- CP-element group 185: 	 branch_block_stmt_271/if_stmt_1062__entry__
      -- CP-element group 185: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/$exit
      -- CP-element group 185: 	 branch_block_stmt_271/if_stmt_1062_dead_link/$entry
      -- CP-element group 185: 	 branch_block_stmt_271/if_stmt_1062_eval_test/$entry
      -- CP-element group 185: 	 branch_block_stmt_271/if_stmt_1062_eval_test/$exit
      -- CP-element group 185: 	 branch_block_stmt_271/if_stmt_1062_eval_test/branch_req
      -- CP-element group 185: 	 branch_block_stmt_271/R_exitcond1_1063_place
      -- CP-element group 185: 	 branch_block_stmt_271/if_stmt_1062_if_link/$entry
      -- CP-element group 185: 	 branch_block_stmt_271/if_stmt_1062_else_link/$entry
      -- 
    branch_req_2328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(185), ack => if_stmt_1062_branch_req_0); -- 
    convTranspose_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_814_elements(179) & convTranspose_CP_814_elements(184);
      gj_convTranspose_cp_element_group_185 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_814_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  merge  transition  place  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	244 
    -- CP-element group 186:  members (13) 
      -- CP-element group 186: 	 branch_block_stmt_271/forx_xend235x_xloopexit_forx_xend235
      -- CP-element group 186: 	 branch_block_stmt_271/merge_stmt_1068__exit__
      -- CP-element group 186: 	 branch_block_stmt_271/if_stmt_1062_if_link/$exit
      -- CP-element group 186: 	 branch_block_stmt_271/if_stmt_1062_if_link/if_choice_transition
      -- CP-element group 186: 	 branch_block_stmt_271/forx_xbody228_forx_xend235x_xloopexit
      -- CP-element group 186: 	 branch_block_stmt_271/forx_xbody228_forx_xend235x_xloopexit_PhiReq/$entry
      -- CP-element group 186: 	 branch_block_stmt_271/forx_xbody228_forx_xend235x_xloopexit_PhiReq/$exit
      -- CP-element group 186: 	 branch_block_stmt_271/merge_stmt_1068_PhiReqMerge
      -- CP-element group 186: 	 branch_block_stmt_271/merge_stmt_1068_PhiAck/$entry
      -- CP-element group 186: 	 branch_block_stmt_271/merge_stmt_1068_PhiAck/$exit
      -- CP-element group 186: 	 branch_block_stmt_271/merge_stmt_1068_PhiAck/dummy
      -- CP-element group 186: 	 branch_block_stmt_271/forx_xend235x_xloopexit_forx_xend235_PhiReq/$entry
      -- CP-element group 186: 	 branch_block_stmt_271/forx_xend235x_xloopexit_forx_xend235_PhiReq/$exit
      -- 
    if_choice_transition_2333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1062_branch_ack_1, ack => convTranspose_CP_814_elements(186)); -- 
    -- CP-element group 187:  fork  transition  place  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	239 
    -- CP-element group 187: 	240 
    -- CP-element group 187:  members (12) 
      -- CP-element group 187: 	 branch_block_stmt_271/forx_xbody228_forx_xbody228
      -- CP-element group 187: 	 branch_block_stmt_271/if_stmt_1062_else_link/$exit
      -- CP-element group 187: 	 branch_block_stmt_271/if_stmt_1062_else_link/else_choice_transition
      -- CP-element group 187: 	 branch_block_stmt_271/forx_xbody228_forx_xbody228_PhiReq/$entry
      -- CP-element group 187: 	 branch_block_stmt_271/forx_xbody228_forx_xbody228_PhiReq/phi_stmt_1031/$entry
      -- CP-element group 187: 	 branch_block_stmt_271/forx_xbody228_forx_xbody228_PhiReq/phi_stmt_1031/phi_stmt_1031_sources/$entry
      -- CP-element group 187: 	 branch_block_stmt_271/forx_xbody228_forx_xbody228_PhiReq/phi_stmt_1031/phi_stmt_1031_sources/type_cast_1037/$entry
      -- CP-element group 187: 	 branch_block_stmt_271/forx_xbody228_forx_xbody228_PhiReq/phi_stmt_1031/phi_stmt_1031_sources/type_cast_1037/SplitProtocol/$entry
      -- CP-element group 187: 	 branch_block_stmt_271/forx_xbody228_forx_xbody228_PhiReq/phi_stmt_1031/phi_stmt_1031_sources/type_cast_1037/SplitProtocol/Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_271/forx_xbody228_forx_xbody228_PhiReq/phi_stmt_1031/phi_stmt_1031_sources/type_cast_1037/SplitProtocol/Sample/rr
      -- CP-element group 187: 	 branch_block_stmt_271/forx_xbody228_forx_xbody228_PhiReq/phi_stmt_1031/phi_stmt_1031_sources/type_cast_1037/SplitProtocol/Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_271/forx_xbody228_forx_xbody228_PhiReq/phi_stmt_1031/phi_stmt_1031_sources/type_cast_1037/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1062_branch_ack_0, ack => convTranspose_CP_814_elements(187)); -- 
    rr_2904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(187), ack => type_cast_1037_inst_req_0); -- 
    cr_2909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(187), ack => type_cast_1037_inst_req_1); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	244 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_271/call_stmt_1072/call_stmt_1072_Sample/cra
      -- CP-element group 188: 	 branch_block_stmt_271/call_stmt_1072/call_stmt_1072_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_271/call_stmt_1072/call_stmt_1072_sample_completed_
      -- 
    cra_2351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1072_call_ack_0, ack => convTranspose_CP_814_elements(188)); -- 
    -- CP-element group 189:  fork  transition  place  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	244 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	247 
    -- CP-element group 189: 	245 
    -- CP-element group 189: 	246 
    -- CP-element group 189:  members (17) 
      -- CP-element group 189: 	 branch_block_stmt_271/call_stmt_1072/call_stmt_1072_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_271/assign_stmt_1079_to_assign_stmt_1095__exit__
      -- CP-element group 189: 	 branch_block_stmt_271/assign_stmt_1079_to_assign_stmt_1095__entry__
      -- CP-element group 189: 	 branch_block_stmt_271/call_stmt_1072__exit__
      -- CP-element group 189: 	 branch_block_stmt_271/forx_xend235_whilex_xbody
      -- CP-element group 189: 	 branch_block_stmt_271/assign_stmt_1079_to_assign_stmt_1095/$entry
      -- CP-element group 189: 	 branch_block_stmt_271/assign_stmt_1079_to_assign_stmt_1095/$exit
      -- CP-element group 189: 	 branch_block_stmt_271/call_stmt_1072/call_stmt_1072_update_completed_
      -- CP-element group 189: 	 branch_block_stmt_271/call_stmt_1072/call_stmt_1072_Update/cca
      -- CP-element group 189: 	 branch_block_stmt_271/call_stmt_1072/$exit
      -- CP-element group 189: 	 branch_block_stmt_271/forx_xend235_whilex_xbody_PhiReq/$entry
      -- CP-element group 189: 	 branch_block_stmt_271/forx_xend235_whilex_xbody_PhiReq/phi_stmt_1098/$entry
      -- CP-element group 189: 	 branch_block_stmt_271/forx_xend235_whilex_xbody_PhiReq/phi_stmt_1098/phi_stmt_1098_sources/$entry
      -- CP-element group 189: 	 branch_block_stmt_271/forx_xend235_whilex_xbody_PhiReq/phi_stmt_1105/$entry
      -- CP-element group 189: 	 branch_block_stmt_271/forx_xend235_whilex_xbody_PhiReq/phi_stmt_1105/phi_stmt_1105_sources/$entry
      -- CP-element group 189: 	 branch_block_stmt_271/forx_xend235_whilex_xbody_PhiReq/phi_stmt_1112/$entry
      -- CP-element group 189: 	 branch_block_stmt_271/forx_xend235_whilex_xbody_PhiReq/phi_stmt_1112/phi_stmt_1112_sources/$entry
      -- 
    cca_2356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1072_call_ack_1, ack => convTranspose_CP_814_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	263 
    -- CP-element group 190: successors 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1182_Sample/ra
      -- CP-element group 190: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1182_Sample/$exit
      -- CP-element group 190: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1182_sample_completed_
      -- 
    ra_2371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1182_inst_ack_0, ack => convTranspose_CP_814_elements(190)); -- 
    -- CP-element group 191:  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	263 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (16) 
      -- CP-element group 191: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_index_computed_1
      -- CP-element group 191: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_index_scaled_1
      -- CP-element group 191: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_index_resize_1/$entry
      -- CP-element group 191: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_index_resize_1/$exit
      -- CP-element group 191: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_index_resize_1/index_resize_req
      -- CP-element group 191: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_index_resize_1/index_resize_ack
      -- CP-element group 191: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_index_scale_1/$entry
      -- CP-element group 191: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_index_scale_1/$exit
      -- CP-element group 191: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_final_index_sum_regn_Sample/req
      -- CP-element group 191: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_final_index_sum_regn_Sample/$entry
      -- CP-element group 191: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_index_resized_1
      -- CP-element group 191: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1182_Update/ca
      -- CP-element group 191: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1182_Update/$exit
      -- CP-element group 191: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1182_update_completed_
      -- CP-element group 191: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_index_scale_1/scale_rename_ack
      -- CP-element group 191: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_index_scale_1/scale_rename_req
      -- 
    ca_2376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1182_inst_ack_1, ack => convTranspose_CP_814_elements(191)); -- 
    req_2401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(191), ack => array_obj_ref_1194_index_offset_req_0); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	211 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_final_index_sum_regn_Sample/ack
      -- CP-element group 192: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_final_index_sum_regn_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_final_index_sum_regn_sample_complete
      -- 
    ack_2402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1194_index_offset_ack_0, ack => convTranspose_CP_814_elements(192)); -- 
    -- CP-element group 193:  transition  input  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	263 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (11) 
      -- CP-element group 193: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1195_request/req
      -- CP-element group 193: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1195_request/$entry
      -- CP-element group 193: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_base_plus_offset/sum_rename_ack
      -- CP-element group 193: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_base_plus_offset/sum_rename_req
      -- CP-element group 193: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_base_plus_offset/$exit
      -- CP-element group 193: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_base_plus_offset/$entry
      -- CP-element group 193: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_final_index_sum_regn_Update/ack
      -- CP-element group 193: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_final_index_sum_regn_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_offset_calculated
      -- CP-element group 193: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_root_address_calculated
      -- CP-element group 193: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1195_sample_start_
      -- 
    ack_2407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1194_index_offset_ack_1, ack => convTranspose_CP_814_elements(193)); -- 
    req_2416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(193), ack => addr_of_1195_final_reg_req_0); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1195_request/$exit
      -- CP-element group 194: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1195_request/ack
      -- CP-element group 194: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1195_sample_completed_
      -- 
    ack_2417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1195_final_reg_ack_0, ack => convTranspose_CP_814_elements(194)); -- 
    -- CP-element group 195:  join  fork  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	263 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (24) 
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1195_complete/$exit
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1195_complete/ack
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_base_address_calculated
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_word_address_calculated
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_root_address_calculated
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_base_address_resized
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_base_addr_resize/$entry
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_base_addr_resize/$exit
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_base_addr_resize/base_resize_req
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_base_addr_resize/base_resize_ack
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_base_plus_offset/$entry
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_base_plus_offset/$exit
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_base_plus_offset/sum_rename_req
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_base_plus_offset/sum_rename_ack
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_word_addrgen/$entry
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_word_addrgen/$exit
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_word_addrgen/root_register_req
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_word_addrgen/root_register_ack
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_Sample/word_access_start/word_0/rr
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_Sample/word_access_start/word_0/$entry
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1195_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_Sample/word_access_start/$entry
      -- CP-element group 195: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_Sample/$entry
      -- 
    ack_2422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1195_final_reg_ack_1, ack => convTranspose_CP_814_elements(195)); -- 
    rr_2455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(195), ack => ptr_deref_1199_load_0_req_0); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (5) 
      -- CP-element group 196: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_Sample/word_access_start/word_0/ra
      -- CP-element group 196: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_Sample/word_access_start/word_0/$exit
      -- CP-element group 196: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_Sample/word_access_start/$exit
      -- CP-element group 196: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_Sample/$exit
      -- 
    ra_2456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1199_load_0_ack_0, ack => convTranspose_CP_814_elements(196)); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	263 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	204 
    -- CP-element group 197:  members (9) 
      -- CP-element group 197: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_Update/word_access_complete/word_0/$exit
      -- CP-element group 197: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_Update/word_access_complete/$exit
      -- CP-element group 197: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_Update/ptr_deref_1199_Merge/merge_ack
      -- CP-element group 197: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_Update/ptr_deref_1199_Merge/merge_req
      -- CP-element group 197: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_Update/ptr_deref_1199_Merge/$exit
      -- CP-element group 197: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_Update/ptr_deref_1199_Merge/$entry
      -- CP-element group 197: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_Update/word_access_complete/word_0/ca
      -- 
    ca_2467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1199_load_0_ack_1, ack => convTranspose_CP_814_elements(197)); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	263 
    -- CP-element group 198: successors 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1203_Sample/ra
      -- CP-element group 198: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1203_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1203_sample_completed_
      -- 
    ra_2481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1203_inst_ack_0, ack => convTranspose_CP_814_elements(198)); -- 
    -- CP-element group 199:  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	263 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (16) 
      -- CP-element group 199: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_final_index_sum_regn_Sample/$entry
      -- CP-element group 199: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_final_index_sum_regn_Sample/req
      -- CP-element group 199: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_index_scale_1/scale_rename_ack
      -- CP-element group 199: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_index_scale_1/scale_rename_req
      -- CP-element group 199: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_index_scale_1/$exit
      -- CP-element group 199: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_index_scale_1/$entry
      -- CP-element group 199: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_index_resize_1/index_resize_ack
      -- CP-element group 199: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_index_resize_1/index_resize_req
      -- CP-element group 199: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_index_resize_1/$exit
      -- CP-element group 199: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_index_resize_1/$entry
      -- CP-element group 199: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_index_computed_1
      -- CP-element group 199: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_index_scaled_1
      -- CP-element group 199: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_index_resized_1
      -- CP-element group 199: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1203_Update/ca
      -- CP-element group 199: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1203_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1203_update_completed_
      -- 
    ca_2486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1203_inst_ack_1, ack => convTranspose_CP_814_elements(199)); -- 
    req_2511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(199), ack => array_obj_ref_1215_index_offset_req_0); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	211 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_final_index_sum_regn_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_final_index_sum_regn_Sample/ack
      -- CP-element group 200: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_final_index_sum_regn_sample_complete
      -- 
    ack_2512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1215_index_offset_ack_0, ack => convTranspose_CP_814_elements(200)); -- 
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	263 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (11) 
      -- CP-element group 201: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_final_index_sum_regn_Update/ack
      -- CP-element group 201: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_final_index_sum_regn_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_base_plus_offset/sum_rename_req
      -- CP-element group 201: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_base_plus_offset/$entry
      -- CP-element group 201: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_base_plus_offset/$exit
      -- CP-element group 201: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_base_plus_offset/sum_rename_ack
      -- CP-element group 201: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1216_request/$entry
      -- CP-element group 201: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1216_request/req
      -- CP-element group 201: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_offset_calculated
      -- CP-element group 201: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_root_address_calculated
      -- CP-element group 201: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1216_sample_start_
      -- 
    ack_2517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1215_index_offset_ack_1, ack => convTranspose_CP_814_elements(201)); -- 
    req_2526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(201), ack => addr_of_1216_final_reg_req_0); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1216_request/$exit
      -- CP-element group 202: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1216_request/ack
      -- CP-element group 202: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1216_sample_completed_
      -- 
    ack_2527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1216_final_reg_ack_0, ack => convTranspose_CP_814_elements(202)); -- 
    -- CP-element group 203:  fork  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	263 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (19) 
      -- CP-element group 203: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1216_complete/$exit
      -- CP-element group 203: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1216_complete/ack
      -- CP-element group 203: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_base_address_calculated
      -- CP-element group 203: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_word_address_calculated
      -- CP-element group 203: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_root_address_calculated
      -- CP-element group 203: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_base_address_resized
      -- CP-element group 203: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_base_addr_resize/$entry
      -- CP-element group 203: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_base_addr_resize/$exit
      -- CP-element group 203: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_base_addr_resize/base_resize_req
      -- CP-element group 203: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1216_update_completed_
      -- CP-element group 203: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_word_addrgen/root_register_ack
      -- CP-element group 203: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_word_addrgen/root_register_req
      -- CP-element group 203: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_word_addrgen/$exit
      -- CP-element group 203: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_word_addrgen/$entry
      -- CP-element group 203: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_base_plus_offset/sum_rename_ack
      -- CP-element group 203: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_base_plus_offset/sum_rename_req
      -- CP-element group 203: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_base_plus_offset/$exit
      -- CP-element group 203: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_base_plus_offset/$entry
      -- CP-element group 203: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_base_addr_resize/base_resize_ack
      -- 
    ack_2532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1216_final_reg_ack_1, ack => convTranspose_CP_814_elements(203)); -- 
    -- CP-element group 204:  join  transition  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	197 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (9) 
      -- CP-element group 204: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_sample_start_
      -- CP-element group 204: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_Sample/word_access_start/word_0/rr
      -- CP-element group 204: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_Sample/word_access_start/word_0/$entry
      -- CP-element group 204: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_Sample/word_access_start/$entry
      -- CP-element group 204: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_Sample/ptr_deref_1219_Split/split_ack
      -- CP-element group 204: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_Sample/ptr_deref_1219_Split/split_req
      -- CP-element group 204: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_Sample/ptr_deref_1219_Split/$exit
      -- CP-element group 204: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_Sample/ptr_deref_1219_Split/$entry
      -- CP-element group 204: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_Sample/$entry
      -- 
    rr_2570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(204), ack => ptr_deref_1219_store_0_req_0); -- 
    convTranspose_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_814_elements(197) & convTranspose_CP_814_elements(203);
      gj_convTranspose_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_814_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (5) 
      -- CP-element group 205: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_Sample/word_access_start/word_0/ra
      -- CP-element group 205: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_Sample/word_access_start/word_0/$exit
      -- CP-element group 205: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_Sample/word_access_start/$exit
      -- CP-element group 205: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_Sample/$exit
      -- 
    ra_2571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1219_store_0_ack_0, ack => convTranspose_CP_814_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	263 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	211 
    -- CP-element group 206:  members (5) 
      -- CP-element group 206: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_Update/word_access_complete/word_0/ca
      -- CP-element group 206: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_Update/word_access_complete/$exit
      -- CP-element group 206: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_Update/word_access_complete/word_0/$exit
      -- CP-element group 206: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_update_completed_
      -- 
    ca_2582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1219_store_0_ack_1, ack => convTranspose_CP_814_elements(206)); -- 
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	263 
    -- CP-element group 207: successors 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1235_sample_completed_
      -- CP-element group 207: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1235_Sample/$exit
      -- CP-element group 207: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1235_Sample/ra
      -- 
    ra_2591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1235_inst_ack_0, ack => convTranspose_CP_814_elements(207)); -- 
    -- CP-element group 208:  transition  input  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	263 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208:  members (6) 
      -- CP-element group 208: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1235_Update/$exit
      -- CP-element group 208: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1235_update_completed_
      -- CP-element group 208: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1256_Sample/rr
      -- CP-element group 208: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1256_Sample/$entry
      -- CP-element group 208: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1256_sample_start_
      -- CP-element group 208: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1235_Update/ca
      -- 
    ca_2596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1235_inst_ack_1, ack => convTranspose_CP_814_elements(208)); -- 
    rr_2604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(208), ack => type_cast_1256_inst_req_0); -- 
    -- CP-element group 209:  transition  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1256_Sample/ra
      -- CP-element group 209: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1256_Sample/$exit
      -- CP-element group 209: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1256_sample_completed_
      -- 
    ra_2605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1256_inst_ack_0, ack => convTranspose_CP_814_elements(209)); -- 
    -- CP-element group 210:  transition  input  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	263 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1256_Update/ca
      -- CP-element group 210: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1256_Update/$exit
      -- CP-element group 210: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1256_update_completed_
      -- 
    ca_2610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1256_inst_ack_1, ack => convTranspose_CP_814_elements(210)); -- 
    -- CP-element group 211:  branch  join  transition  place  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	206 
    -- CP-element group 211: 	192 
    -- CP-element group 211: 	200 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	212 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (10) 
      -- CP-element group 211: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274__exit__
      -- CP-element group 211: 	 branch_block_stmt_271/if_stmt_1275__entry__
      -- CP-element group 211: 	 branch_block_stmt_271/if_stmt_1275_else_link/$entry
      -- CP-element group 211: 	 branch_block_stmt_271/if_stmt_1275_if_link/$entry
      -- CP-element group 211: 	 branch_block_stmt_271/if_stmt_1275_eval_test/branch_req
      -- CP-element group 211: 	 branch_block_stmt_271/if_stmt_1275_eval_test/$exit
      -- CP-element group 211: 	 branch_block_stmt_271/if_stmt_1275_eval_test/$entry
      -- CP-element group 211: 	 branch_block_stmt_271/if_stmt_1275_dead_link/$entry
      -- CP-element group 211: 	 branch_block_stmt_271/R_cmp342_1276_place
      -- CP-element group 211: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/$exit
      -- 
    branch_req_2618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(211), ack => if_stmt_1275_branch_req_0); -- 
    convTranspose_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTranspose_CP_814_elements(206) & convTranspose_CP_814_elements(192) & convTranspose_CP_814_elements(200) & convTranspose_CP_814_elements(210);
      gj_convTranspose_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_814_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	211 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	214 
    -- CP-element group 212: 	215 
    -- CP-element group 212:  members (18) 
      -- CP-element group 212: 	 branch_block_stmt_271/assign_stmt_1287__entry__
      -- CP-element group 212: 	 branch_block_stmt_271/merge_stmt_1281__exit__
      -- CP-element group 212: 	 branch_block_stmt_271/assign_stmt_1287/type_cast_1286_Update/cr
      -- CP-element group 212: 	 branch_block_stmt_271/assign_stmt_1287/type_cast_1286_Update/$entry
      -- CP-element group 212: 	 branch_block_stmt_271/assign_stmt_1287/type_cast_1286_Sample/rr
      -- CP-element group 212: 	 branch_block_stmt_271/assign_stmt_1287/type_cast_1286_Sample/$entry
      -- CP-element group 212: 	 branch_block_stmt_271/assign_stmt_1287/type_cast_1286_update_start_
      -- CP-element group 212: 	 branch_block_stmt_271/assign_stmt_1287/type_cast_1286_sample_start_
      -- CP-element group 212: 	 branch_block_stmt_271/assign_stmt_1287/$entry
      -- CP-element group 212: 	 branch_block_stmt_271/if_stmt_1275_if_link/if_choice_transition
      -- CP-element group 212: 	 branch_block_stmt_271/if_stmt_1275_if_link/$exit
      -- CP-element group 212: 	 branch_block_stmt_271/whilex_xbody_whilex_xend
      -- CP-element group 212: 	 branch_block_stmt_271/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 212: 	 branch_block_stmt_271/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 212: 	 branch_block_stmt_271/merge_stmt_1281_PhiReqMerge
      -- CP-element group 212: 	 branch_block_stmt_271/merge_stmt_1281_PhiAck/$entry
      -- CP-element group 212: 	 branch_block_stmt_271/merge_stmt_1281_PhiAck/$exit
      -- CP-element group 212: 	 branch_block_stmt_271/merge_stmt_1281_PhiAck/dummy
      -- 
    if_choice_transition_2623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1275_branch_ack_1, ack => convTranspose_CP_814_elements(212)); -- 
    cr_2645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(212), ack => type_cast_1286_inst_req_1); -- 
    rr_2640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(212), ack => type_cast_1286_inst_req_0); -- 
    -- CP-element group 213:  fork  transition  place  input  output  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	249 
    -- CP-element group 213: 	250 
    -- CP-element group 213: 	256 
    -- CP-element group 213: 	252 
    -- CP-element group 213: 	253 
    -- CP-element group 213: 	255 
    -- CP-element group 213:  members (28) 
      -- CP-element group 213: 	 branch_block_stmt_271/if_stmt_1275_else_link/else_choice_transition
      -- CP-element group 213: 	 branch_block_stmt_271/if_stmt_1275_else_link/$exit
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/$entry
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1098/$entry
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1098/phi_stmt_1098_sources/$entry
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1098/phi_stmt_1098_sources/type_cast_1104/$entry
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1098/phi_stmt_1098_sources/type_cast_1104/SplitProtocol/$entry
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1098/phi_stmt_1098_sources/type_cast_1104/SplitProtocol/Sample/$entry
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1098/phi_stmt_1098_sources/type_cast_1104/SplitProtocol/Sample/rr
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1098/phi_stmt_1098_sources/type_cast_1104/SplitProtocol/Update/$entry
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1098/phi_stmt_1098_sources/type_cast_1104/SplitProtocol/Update/cr
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1105/$entry
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1105/phi_stmt_1105_sources/$entry
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1105/phi_stmt_1105_sources/type_cast_1111/$entry
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1105/phi_stmt_1105_sources/type_cast_1111/SplitProtocol/$entry
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1105/phi_stmt_1105_sources/type_cast_1111/SplitProtocol/Sample/$entry
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1105/phi_stmt_1105_sources/type_cast_1111/SplitProtocol/Sample/rr
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1105/phi_stmt_1105_sources/type_cast_1111/SplitProtocol/Update/$entry
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1105/phi_stmt_1105_sources/type_cast_1111/SplitProtocol/Update/cr
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1112/$entry
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1112/phi_stmt_1112_sources/$entry
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1112/phi_stmt_1112_sources/type_cast_1118/$entry
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1112/phi_stmt_1112_sources/type_cast_1118/SplitProtocol/$entry
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1112/phi_stmt_1112_sources/type_cast_1118/SplitProtocol/Sample/$entry
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1112/phi_stmt_1112_sources/type_cast_1118/SplitProtocol/Sample/rr
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1112/phi_stmt_1112_sources/type_cast_1118/SplitProtocol/Update/$entry
      -- CP-element group 213: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1112/phi_stmt_1112_sources/type_cast_1118/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1275_branch_ack_0, ack => convTranspose_CP_814_elements(213)); -- 
    rr_2985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(213), ack => type_cast_1104_inst_req_0); -- 
    cr_2990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(213), ack => type_cast_1104_inst_req_1); -- 
    rr_3008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(213), ack => type_cast_1111_inst_req_0); -- 
    cr_3013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(213), ack => type_cast_1111_inst_req_1); -- 
    rr_3031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(213), ack => type_cast_1118_inst_req_0); -- 
    cr_3036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(213), ack => type_cast_1118_inst_req_1); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	212 
    -- CP-element group 214: successors 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_271/assign_stmt_1287/type_cast_1286_Sample/ra
      -- CP-element group 214: 	 branch_block_stmt_271/assign_stmt_1287/type_cast_1286_Sample/$exit
      -- CP-element group 214: 	 branch_block_stmt_271/assign_stmt_1287/type_cast_1286_sample_completed_
      -- 
    ra_2641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1286_inst_ack_0, ack => convTranspose_CP_814_elements(214)); -- 
    -- CP-element group 215:  fork  transition  place  input  output  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	212 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215: 	217 
    -- CP-element group 215: 	219 
    -- CP-element group 215:  members (16) 
      -- CP-element group 215: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/call_stmt_1290_sample_start_
      -- CP-element group 215: 	 branch_block_stmt_271/assign_stmt_1287__exit__
      -- CP-element group 215: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303__entry__
      -- CP-element group 215: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/call_stmt_1290_update_start_
      -- CP-element group 215: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/type_cast_1294_Update/$entry
      -- CP-element group 215: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/call_stmt_1290_Sample/$entry
      -- CP-element group 215: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/call_stmt_1290_Sample/crr
      -- CP-element group 215: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/call_stmt_1290_Update/$entry
      -- CP-element group 215: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/call_stmt_1290_Update/ccr
      -- CP-element group 215: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/type_cast_1294_update_start_
      -- CP-element group 215: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/$entry
      -- CP-element group 215: 	 branch_block_stmt_271/assign_stmt_1287/type_cast_1286_Update/ca
      -- CP-element group 215: 	 branch_block_stmt_271/assign_stmt_1287/type_cast_1286_Update/$exit
      -- CP-element group 215: 	 branch_block_stmt_271/assign_stmt_1287/type_cast_1286_update_completed_
      -- CP-element group 215: 	 branch_block_stmt_271/assign_stmt_1287/$exit
      -- CP-element group 215: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/type_cast_1294_Update/cr
      -- 
    ca_2646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1286_inst_ack_1, ack => convTranspose_CP_814_elements(215)); -- 
    crr_2657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(215), ack => call_stmt_1290_call_req_0); -- 
    ccr_2662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(215), ack => call_stmt_1290_call_req_1); -- 
    cr_2676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(215), ack => type_cast_1294_inst_req_1); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/call_stmt_1290_sample_completed_
      -- CP-element group 216: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/call_stmt_1290_Sample/$exit
      -- CP-element group 216: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/call_stmt_1290_Sample/cra
      -- 
    cra_2658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1290_call_ack_0, ack => convTranspose_CP_814_elements(216)); -- 
    -- CP-element group 217:  transition  input  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	215 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (6) 
      -- CP-element group 217: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/call_stmt_1290_update_completed_
      -- CP-element group 217: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/call_stmt_1290_Update/$exit
      -- CP-element group 217: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/call_stmt_1290_Update/cca
      -- CP-element group 217: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/type_cast_1294_sample_start_
      -- CP-element group 217: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/type_cast_1294_Sample/$entry
      -- CP-element group 217: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/type_cast_1294_Sample/rr
      -- 
    cca_2663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1290_call_ack_1, ack => convTranspose_CP_814_elements(217)); -- 
    rr_2671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(217), ack => type_cast_1294_inst_req_0); -- 
    -- CP-element group 218:  transition  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/type_cast_1294_sample_completed_
      -- CP-element group 218: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/type_cast_1294_Sample/$exit
      -- CP-element group 218: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/type_cast_1294_Sample/ra
      -- 
    ra_2672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1294_inst_ack_0, ack => convTranspose_CP_814_elements(218)); -- 
    -- CP-element group 219:  transition  input  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	215 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	220 
    -- CP-element group 219:  members (6) 
      -- CP-element group 219: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/type_cast_1294_update_completed_
      -- CP-element group 219: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/WPIPE_elapsed_time_pipe_1301_Sample/req
      -- CP-element group 219: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/WPIPE_elapsed_time_pipe_1301_Sample/$entry
      -- CP-element group 219: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/WPIPE_elapsed_time_pipe_1301_sample_start_
      -- CP-element group 219: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/type_cast_1294_Update/ca
      -- CP-element group 219: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/type_cast_1294_Update/$exit
      -- 
    ca_2677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1294_inst_ack_1, ack => convTranspose_CP_814_elements(219)); -- 
    req_2685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(219), ack => WPIPE_elapsed_time_pipe_1301_inst_req_0); -- 
    -- CP-element group 220:  transition  input  output  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	219 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	221 
    -- CP-element group 220:  members (6) 
      -- CP-element group 220: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/WPIPE_elapsed_time_pipe_1301_Update/req
      -- CP-element group 220: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/WPIPE_elapsed_time_pipe_1301_Update/$entry
      -- CP-element group 220: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/WPIPE_elapsed_time_pipe_1301_Sample/ack
      -- CP-element group 220: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/WPIPE_elapsed_time_pipe_1301_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/WPIPE_elapsed_time_pipe_1301_update_start_
      -- CP-element group 220: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/WPIPE_elapsed_time_pipe_1301_sample_completed_
      -- 
    ack_2686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1301_inst_ack_0, ack => convTranspose_CP_814_elements(220)); -- 
    req_2690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(220), ack => WPIPE_elapsed_time_pipe_1301_inst_req_1); -- 
    -- CP-element group 221:  fork  transition  place  input  output  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	220 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	222 
    -- CP-element group 221: 	223 
    -- CP-element group 221:  members (13) 
      -- CP-element group 221: 	 branch_block_stmt_271/call_stmt_1306__entry__
      -- CP-element group 221: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303__exit__
      -- CP-element group 221: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/$exit
      -- CP-element group 221: 	 branch_block_stmt_271/call_stmt_1306/call_stmt_1306_Update/ccr
      -- CP-element group 221: 	 branch_block_stmt_271/call_stmt_1306/call_stmt_1306_Update/$entry
      -- CP-element group 221: 	 branch_block_stmt_271/call_stmt_1306/$entry
      -- CP-element group 221: 	 branch_block_stmt_271/call_stmt_1306/call_stmt_1306_Sample/crr
      -- CP-element group 221: 	 branch_block_stmt_271/call_stmt_1306/call_stmt_1306_Sample/$entry
      -- CP-element group 221: 	 branch_block_stmt_271/call_stmt_1306/call_stmt_1306_update_start_
      -- CP-element group 221: 	 branch_block_stmt_271/call_stmt_1306/call_stmt_1306_sample_start_
      -- CP-element group 221: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/WPIPE_elapsed_time_pipe_1301_Update/ack
      -- CP-element group 221: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/WPIPE_elapsed_time_pipe_1301_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_271/call_stmt_1290_to_assign_stmt_1303/WPIPE_elapsed_time_pipe_1301_update_completed_
      -- 
    ack_2691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1301_inst_ack_1, ack => convTranspose_CP_814_elements(221)); -- 
    ccr_2707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(221), ack => call_stmt_1306_call_req_1); -- 
    crr_2702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(221), ack => call_stmt_1306_call_req_0); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	221 
    -- CP-element group 222: successors 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_271/call_stmt_1306/call_stmt_1306_Sample/cra
      -- CP-element group 222: 	 branch_block_stmt_271/call_stmt_1306/call_stmt_1306_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_271/call_stmt_1306/call_stmt_1306_sample_completed_
      -- 
    cra_2703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1306_call_ack_0, ack => convTranspose_CP_814_elements(222)); -- 
    -- CP-element group 223:  transition  place  input  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	221 
    -- CP-element group 223: successors 
    -- CP-element group 223:  members (16) 
      -- CP-element group 223: 	 $exit
      -- CP-element group 223: 	 branch_block_stmt_271/branch_block_stmt_271__exit__
      -- CP-element group 223: 	 branch_block_stmt_271/$exit
      -- CP-element group 223: 	 branch_block_stmt_271/merge_stmt_1308__exit__
      -- CP-element group 223: 	 branch_block_stmt_271/return__
      -- CP-element group 223: 	 branch_block_stmt_271/call_stmt_1306__exit__
      -- CP-element group 223: 	 branch_block_stmt_271/call_stmt_1306/call_stmt_1306_Update/cca
      -- CP-element group 223: 	 branch_block_stmt_271/call_stmt_1306/call_stmt_1306_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_271/call_stmt_1306/call_stmt_1306_update_completed_
      -- CP-element group 223: 	 branch_block_stmt_271/call_stmt_1306/$exit
      -- CP-element group 223: 	 branch_block_stmt_271/return___PhiReq/$entry
      -- CP-element group 223: 	 branch_block_stmt_271/return___PhiReq/$exit
      -- CP-element group 223: 	 branch_block_stmt_271/merge_stmt_1308_PhiReqMerge
      -- CP-element group 223: 	 branch_block_stmt_271/merge_stmt_1308_PhiAck/$entry
      -- CP-element group 223: 	 branch_block_stmt_271/merge_stmt_1308_PhiAck/$exit
      -- CP-element group 223: 	 branch_block_stmt_271/merge_stmt_1308_PhiAck/dummy
      -- 
    cca_2708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1306_call_ack_1, ack => convTranspose_CP_814_elements(223)); -- 
    -- CP-element group 224:  transition  output  delay-element  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	124 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	228 
    -- CP-element group 224:  members (5) 
      -- CP-element group 224: 	 branch_block_stmt_271/bbx_xnph378_forx_xbody_PhiReq/$exit
      -- CP-element group 224: 	 branch_block_stmt_271/bbx_xnph378_forx_xbody_PhiReq/phi_stmt_712/$exit
      -- CP-element group 224: 	 branch_block_stmt_271/bbx_xnph378_forx_xbody_PhiReq/phi_stmt_712/phi_stmt_712_req
      -- CP-element group 224: 	 branch_block_stmt_271/bbx_xnph378_forx_xbody_PhiReq/phi_stmt_712/phi_stmt_712_sources/type_cast_716_konst_delay_trans
      -- CP-element group 224: 	 branch_block_stmt_271/bbx_xnph378_forx_xbody_PhiReq/phi_stmt_712/phi_stmt_712_sources/$exit
      -- 
    phi_stmt_712_req_2731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_712_req_2731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(224), ack => phi_stmt_712_req_0); -- 
    -- Element group convTranspose_CP_814_elements(224) is a control-delay.
    cp_element_224_delay: control_delay_element  generic map(name => " 224_delay", delay_value => 1)  port map(req => convTranspose_CP_814_elements(124), ack => convTranspose_CP_814_elements(224), clk => clk, reset =>reset);
    -- CP-element group 225:  transition  input  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	166 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	227 
    -- CP-element group 225:  members (2) 
      -- CP-element group 225: 	 branch_block_stmt_271/forx_xbody_forx_xbody_PhiReq/phi_stmt_712/phi_stmt_712_sources/type_cast_718/SplitProtocol/Sample/ra
      -- CP-element group 225: 	 branch_block_stmt_271/forx_xbody_forx_xbody_PhiReq/phi_stmt_712/phi_stmt_712_sources/type_cast_718/SplitProtocol/Sample/$exit
      -- 
    ra_2751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_718_inst_ack_0, ack => convTranspose_CP_814_elements(225)); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	166 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	227 
    -- CP-element group 226:  members (2) 
      -- CP-element group 226: 	 branch_block_stmt_271/forx_xbody_forx_xbody_PhiReq/phi_stmt_712/phi_stmt_712_sources/type_cast_718/SplitProtocol/Update/ca
      -- CP-element group 226: 	 branch_block_stmt_271/forx_xbody_forx_xbody_PhiReq/phi_stmt_712/phi_stmt_712_sources/type_cast_718/SplitProtocol/Update/$exit
      -- 
    ca_2756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_718_inst_ack_1, ack => convTranspose_CP_814_elements(226)); -- 
    -- CP-element group 227:  join  transition  output  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	225 
    -- CP-element group 227: 	226 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (6) 
      -- CP-element group 227: 	 branch_block_stmt_271/forx_xbody_forx_xbody_PhiReq/phi_stmt_712/phi_stmt_712_req
      -- CP-element group 227: 	 branch_block_stmt_271/forx_xbody_forx_xbody_PhiReq/phi_stmt_712/phi_stmt_712_sources/type_cast_718/SplitProtocol/$exit
      -- CP-element group 227: 	 branch_block_stmt_271/forx_xbody_forx_xbody_PhiReq/phi_stmt_712/phi_stmt_712_sources/type_cast_718/$exit
      -- CP-element group 227: 	 branch_block_stmt_271/forx_xbody_forx_xbody_PhiReq/phi_stmt_712/phi_stmt_712_sources/$exit
      -- CP-element group 227: 	 branch_block_stmt_271/forx_xbody_forx_xbody_PhiReq/phi_stmt_712/$exit
      -- CP-element group 227: 	 branch_block_stmt_271/forx_xbody_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_712_req_2757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_712_req_2757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(227), ack => phi_stmt_712_req_1); -- 
    convTranspose_cp_element_group_227: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_227"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_814_elements(225) & convTranspose_CP_814_elements(226);
      gj_convTranspose_cp_element_group_227 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_814_elements(227), clk => clk, reset => reset); --
    end block;
    -- CP-element group 228:  merge  transition  place  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	227 
    -- CP-element group 228: 	224 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228:  members (2) 
      -- CP-element group 228: 	 branch_block_stmt_271/merge_stmt_711_PhiReqMerge
      -- CP-element group 228: 	 branch_block_stmt_271/merge_stmt_711_PhiAck/$entry
      -- 
    convTranspose_CP_814_elements(228) <= OrReduce(convTranspose_CP_814_elements(227) & convTranspose_CP_814_elements(224));
    -- CP-element group 229:  fork  transition  place  input  output  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	148 
    -- CP-element group 229: 	152 
    -- CP-element group 229: 	156 
    -- CP-element group 229: 	160 
    -- CP-element group 229: 	129 
    -- CP-element group 229: 	132 
    -- CP-element group 229: 	163 
    -- CP-element group 229: 	125 
    -- CP-element group 229: 	126 
    -- CP-element group 229: 	128 
    -- CP-element group 229: 	144 
    -- CP-element group 229: 	140 
    -- CP-element group 229: 	136 
    -- CP-element group 229:  members (56) 
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_728_Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/$entry
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_728_Sample/rr
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_index_resize_1/index_resize_ack
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/addr_of_725_complete/$entry
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/addr_of_725_complete/req
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_index_resize_1/$entry
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_index_computed_1
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_index_resize_1/$exit
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_745_Update/cr
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/RPIPE_ConvTranspose_input_pipe_728_sample_start_
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_index_scaled_1
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_index_scale_1/$entry
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_index_scale_1/$exit
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_index_scale_1/scale_rename_req
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_index_scale_1/scale_rename_ack
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_732_update_start_
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_index_resize_1/index_resize_req
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874__entry__
      -- CP-element group 229: 	 branch_block_stmt_271/merge_stmt_711__exit__
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_final_index_sum_regn_update_start
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_final_index_sum_regn_Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_745_update_start_
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_index_resized_1
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_final_index_sum_regn_Update/req
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_745_Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_final_index_sum_regn_Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/array_obj_ref_724_final_index_sum_regn_Sample/req
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_732_Update/cr
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_732_Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/addr_of_725_update_start_
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_763_update_start_
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_763_Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_763_Update/cr
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_781_update_start_
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_781_Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_781_Update/cr
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_799_update_start_
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_799_Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_799_Update/cr
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_817_update_start_
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_817_Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_817_Update/cr
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_835_update_start_
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_835_Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_835_Update/cr
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_853_update_start_
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_853_Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/type_cast_853_Update/cr
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_update_start_
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_Update/word_access_complete/$entry
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_Update/word_access_complete/word_0/$entry
      -- CP-element group 229: 	 branch_block_stmt_271/assign_stmt_726_to_assign_stmt_874/ptr_deref_861_Update/word_access_complete/word_0/cr
      -- CP-element group 229: 	 branch_block_stmt_271/merge_stmt_711_PhiAck/phi_stmt_712_ack
      -- CP-element group 229: 	 branch_block_stmt_271/merge_stmt_711_PhiAck/$exit
      -- 
    phi_stmt_712_ack_2762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_712_ack_0, ack => convTranspose_CP_814_elements(229)); -- 
    rr_1822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(229), ack => RPIPE_ConvTranspose_input_pipe_728_inst_req_0); -- 
    req_1813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(229), ack => addr_of_725_final_reg_req_1); -- 
    cr_1869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(229), ack => type_cast_745_inst_req_1); -- 
    req_1798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(229), ack => array_obj_ref_724_index_offset_req_1); -- 
    req_1793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(229), ack => array_obj_ref_724_index_offset_req_0); -- 
    cr_1841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(229), ack => type_cast_732_inst_req_1); -- 
    cr_1897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(229), ack => type_cast_763_inst_req_1); -- 
    cr_1925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(229), ack => type_cast_781_inst_req_1); -- 
    cr_1953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(229), ack => type_cast_799_inst_req_1); -- 
    cr_1981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(229), ack => type_cast_817_inst_req_1); -- 
    cr_2009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(229), ack => type_cast_835_inst_req_1); -- 
    cr_2037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(229), ack => type_cast_853_inst_req_1); -- 
    cr_2087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(229), ack => ptr_deref_861_store_0_req_1); -- 
    -- CP-element group 230:  merge  branch  transition  place  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	122 
    -- CP-element group 230: 	165 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	167 
    -- CP-element group 230: 	168 
    -- CP-element group 230:  members (17) 
      -- CP-element group 230: 	 branch_block_stmt_271/if_stmt_891__entry__
      -- CP-element group 230: 	 branch_block_stmt_271/assign_stmt_890__exit__
      -- CP-element group 230: 	 branch_block_stmt_271/merge_stmt_883_PhiAck/$exit
      -- CP-element group 230: 	 branch_block_stmt_271/merge_stmt_883_PhiAck/dummy
      -- CP-element group 230: 	 branch_block_stmt_271/assign_stmt_890__entry__
      -- CP-element group 230: 	 branch_block_stmt_271/merge_stmt_883__exit__
      -- CP-element group 230: 	 branch_block_stmt_271/merge_stmt_883_PhiAck/$entry
      -- CP-element group 230: 	 branch_block_stmt_271/merge_stmt_883_PhiReqMerge
      -- CP-element group 230: 	 branch_block_stmt_271/assign_stmt_890/$entry
      -- CP-element group 230: 	 branch_block_stmt_271/assign_stmt_890/$exit
      -- CP-element group 230: 	 branch_block_stmt_271/if_stmt_891_dead_link/$entry
      -- CP-element group 230: 	 branch_block_stmt_271/if_stmt_891_eval_test/$entry
      -- CP-element group 230: 	 branch_block_stmt_271/if_stmt_891_eval_test/$exit
      -- CP-element group 230: 	 branch_block_stmt_271/if_stmt_891_eval_test/branch_req
      -- CP-element group 230: 	 branch_block_stmt_271/R_cmp212372_892_place
      -- CP-element group 230: 	 branch_block_stmt_271/if_stmt_891_if_link/$entry
      -- CP-element group 230: 	 branch_block_stmt_271/if_stmt_891_else_link/$entry
      -- 
    branch_req_2118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(230), ack => if_stmt_891_branch_req_0); -- 
    convTranspose_CP_814_elements(230) <= OrReduce(convTranspose_CP_814_elements(122) & convTranspose_CP_814_elements(165));
    -- CP-element group 231:  transition  output  delay-element  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	170 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	235 
    -- CP-element group 231:  members (5) 
      -- CP-element group 231: 	 branch_block_stmt_271/bbx_xnph374_forx_xbody214_PhiReq/phi_stmt_950/phi_stmt_950_sources/$exit
      -- CP-element group 231: 	 branch_block_stmt_271/bbx_xnph374_forx_xbody214_PhiReq/phi_stmt_950/phi_stmt_950_sources/type_cast_954_konst_delay_trans
      -- CP-element group 231: 	 branch_block_stmt_271/bbx_xnph374_forx_xbody214_PhiReq/phi_stmt_950/phi_stmt_950_req
      -- CP-element group 231: 	 branch_block_stmt_271/bbx_xnph374_forx_xbody214_PhiReq/phi_stmt_950/$exit
      -- CP-element group 231: 	 branch_block_stmt_271/bbx_xnph374_forx_xbody214_PhiReq/$exit
      -- 
    phi_stmt_950_req_2808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_950_req_2808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(231), ack => phi_stmt_950_req_0); -- 
    -- Element group convTranspose_CP_814_elements(231) is a control-delay.
    cp_element_231_delay: control_delay_element  generic map(name => " 231_delay", delay_value => 1)  port map(req => convTranspose_CP_814_elements(170), ack => convTranspose_CP_814_elements(231), clk => clk, reset =>reset);
    -- CP-element group 232:  transition  input  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	174 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	234 
    -- CP-element group 232:  members (2) 
      -- CP-element group 232: 	 branch_block_stmt_271/forx_xbody214_forx_xbody214_PhiReq/phi_stmt_950/phi_stmt_950_sources/type_cast_956/SplitProtocol/Sample/$exit
      -- CP-element group 232: 	 branch_block_stmt_271/forx_xbody214_forx_xbody214_PhiReq/phi_stmt_950/phi_stmt_950_sources/type_cast_956/SplitProtocol/Sample/ra
      -- 
    ra_2828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_956_inst_ack_0, ack => convTranspose_CP_814_elements(232)); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	174 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	234 
    -- CP-element group 233:  members (2) 
      -- CP-element group 233: 	 branch_block_stmt_271/forx_xbody214_forx_xbody214_PhiReq/phi_stmt_950/phi_stmt_950_sources/type_cast_956/SplitProtocol/Update/ca
      -- CP-element group 233: 	 branch_block_stmt_271/forx_xbody214_forx_xbody214_PhiReq/phi_stmt_950/phi_stmt_950_sources/type_cast_956/SplitProtocol/Update/$exit
      -- 
    ca_2833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_956_inst_ack_1, ack => convTranspose_CP_814_elements(233)); -- 
    -- CP-element group 234:  join  transition  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	232 
    -- CP-element group 234: 	233 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234:  members (6) 
      -- CP-element group 234: 	 branch_block_stmt_271/forx_xbody214_forx_xbody214_PhiReq/phi_stmt_950/phi_stmt_950_req
      -- CP-element group 234: 	 branch_block_stmt_271/forx_xbody214_forx_xbody214_PhiReq/phi_stmt_950/phi_stmt_950_sources/type_cast_956/SplitProtocol/$exit
      -- CP-element group 234: 	 branch_block_stmt_271/forx_xbody214_forx_xbody214_PhiReq/phi_stmt_950/phi_stmt_950_sources/type_cast_956/$exit
      -- CP-element group 234: 	 branch_block_stmt_271/forx_xbody214_forx_xbody214_PhiReq/phi_stmt_950/phi_stmt_950_sources/$exit
      -- CP-element group 234: 	 branch_block_stmt_271/forx_xbody214_forx_xbody214_PhiReq/phi_stmt_950/$exit
      -- CP-element group 234: 	 branch_block_stmt_271/forx_xbody214_forx_xbody214_PhiReq/$exit
      -- 
    phi_stmt_950_req_2834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_950_req_2834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(234), ack => phi_stmt_950_req_1); -- 
    convTranspose_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_814_elements(232) & convTranspose_CP_814_elements(233);
      gj_convTranspose_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_814_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  merge  transition  place  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	231 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (2) 
      -- CP-element group 235: 	 branch_block_stmt_271/merge_stmt_949_PhiAck/$entry
      -- CP-element group 235: 	 branch_block_stmt_271/merge_stmt_949_PhiReqMerge
      -- 
    convTranspose_CP_814_elements(235) <= OrReduce(convTranspose_CP_814_elements(231) & convTranspose_CP_814_elements(234));
    -- CP-element group 236:  fork  transition  place  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	171 
    -- CP-element group 236: 	172 
    -- CP-element group 236:  members (11) 
      -- CP-element group 236: 	 branch_block_stmt_271/merge_stmt_949__exit__
      -- CP-element group 236: 	 branch_block_stmt_271/call_stmt_959_to_assign_stmt_970__entry__
      -- CP-element group 236: 	 branch_block_stmt_271/merge_stmt_949_PhiAck/phi_stmt_950_ack
      -- CP-element group 236: 	 branch_block_stmt_271/merge_stmt_949_PhiAck/$exit
      -- CP-element group 236: 	 branch_block_stmt_271/call_stmt_959_to_assign_stmt_970/$entry
      -- CP-element group 236: 	 branch_block_stmt_271/call_stmt_959_to_assign_stmt_970/call_stmt_959_sample_start_
      -- CP-element group 236: 	 branch_block_stmt_271/call_stmt_959_to_assign_stmt_970/call_stmt_959_update_start_
      -- CP-element group 236: 	 branch_block_stmt_271/call_stmt_959_to_assign_stmt_970/call_stmt_959_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_271/call_stmt_959_to_assign_stmt_970/call_stmt_959_Sample/crr
      -- CP-element group 236: 	 branch_block_stmt_271/call_stmt_959_to_assign_stmt_970/call_stmt_959_Update/$entry
      -- CP-element group 236: 	 branch_block_stmt_271/call_stmt_959_to_assign_stmt_970/call_stmt_959_Update/ccr
      -- 
    phi_stmt_950_ack_2839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_950_ack_0, ack => convTranspose_CP_814_elements(236)); -- 
    crr_2157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(236), ack => call_stmt_959_call_req_0); -- 
    ccr_2162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(236), ack => call_stmt_959_call_req_1); -- 
    -- CP-element group 237:  merge  branch  transition  place  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	168 
    -- CP-element group 237: 	173 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	175 
    -- CP-element group 237: 	176 
    -- CP-element group 237:  members (17) 
      -- CP-element group 237: 	 branch_block_stmt_271/if_stmt_987__entry__
      -- CP-element group 237: 	 branch_block_stmt_271/assign_stmt_986__exit__
      -- CP-element group 237: 	 branch_block_stmt_271/assign_stmt_986__entry__
      -- CP-element group 237: 	 branch_block_stmt_271/merge_stmt_979__exit__
      -- CP-element group 237: 	 branch_block_stmt_271/assign_stmt_986/$entry
      -- CP-element group 237: 	 branch_block_stmt_271/assign_stmt_986/$exit
      -- CP-element group 237: 	 branch_block_stmt_271/if_stmt_987_dead_link/$entry
      -- CP-element group 237: 	 branch_block_stmt_271/if_stmt_987_eval_test/$entry
      -- CP-element group 237: 	 branch_block_stmt_271/if_stmt_987_eval_test/$exit
      -- CP-element group 237: 	 branch_block_stmt_271/if_stmt_987_eval_test/branch_req
      -- CP-element group 237: 	 branch_block_stmt_271/R_cmp226369_988_place
      -- CP-element group 237: 	 branch_block_stmt_271/if_stmt_987_if_link/$entry
      -- CP-element group 237: 	 branch_block_stmt_271/if_stmt_987_else_link/$entry
      -- CP-element group 237: 	 branch_block_stmt_271/merge_stmt_979_PhiReqMerge
      -- CP-element group 237: 	 branch_block_stmt_271/merge_stmt_979_PhiAck/$entry
      -- CP-element group 237: 	 branch_block_stmt_271/merge_stmt_979_PhiAck/$exit
      -- CP-element group 237: 	 branch_block_stmt_271/merge_stmt_979_PhiAck/dummy
      -- 
    branch_req_2193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(237), ack => if_stmt_987_branch_req_0); -- 
    convTranspose_CP_814_elements(237) <= OrReduce(convTranspose_CP_814_elements(168) & convTranspose_CP_814_elements(173));
    -- CP-element group 238:  transition  output  delay-element  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	178 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	242 
    -- CP-element group 238:  members (5) 
      -- CP-element group 238: 	 branch_block_stmt_271/bbx_xnph_forx_xbody228_PhiReq/$exit
      -- CP-element group 238: 	 branch_block_stmt_271/bbx_xnph_forx_xbody228_PhiReq/phi_stmt_1031/$exit
      -- CP-element group 238: 	 branch_block_stmt_271/bbx_xnph_forx_xbody228_PhiReq/phi_stmt_1031/phi_stmt_1031_sources/$exit
      -- CP-element group 238: 	 branch_block_stmt_271/bbx_xnph_forx_xbody228_PhiReq/phi_stmt_1031/phi_stmt_1031_sources/type_cast_1035_konst_delay_trans
      -- CP-element group 238: 	 branch_block_stmt_271/bbx_xnph_forx_xbody228_PhiReq/phi_stmt_1031/phi_stmt_1031_req
      -- 
    phi_stmt_1031_req_2885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1031_req_2885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(238), ack => phi_stmt_1031_req_0); -- 
    -- Element group convTranspose_CP_814_elements(238) is a control-delay.
    cp_element_238_delay: control_delay_element  generic map(name => " 238_delay", delay_value => 1)  port map(req => convTranspose_CP_814_elements(178), ack => convTranspose_CP_814_elements(238), clk => clk, reset =>reset);
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	187 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	241 
    -- CP-element group 239:  members (2) 
      -- CP-element group 239: 	 branch_block_stmt_271/forx_xbody228_forx_xbody228_PhiReq/phi_stmt_1031/phi_stmt_1031_sources/type_cast_1037/SplitProtocol/Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_271/forx_xbody228_forx_xbody228_PhiReq/phi_stmt_1031/phi_stmt_1031_sources/type_cast_1037/SplitProtocol/Sample/ra
      -- 
    ra_2905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1037_inst_ack_0, ack => convTranspose_CP_814_elements(239)); -- 
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	187 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (2) 
      -- CP-element group 240: 	 branch_block_stmt_271/forx_xbody228_forx_xbody228_PhiReq/phi_stmt_1031/phi_stmt_1031_sources/type_cast_1037/SplitProtocol/Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_271/forx_xbody228_forx_xbody228_PhiReq/phi_stmt_1031/phi_stmt_1031_sources/type_cast_1037/SplitProtocol/Update/ca
      -- 
    ca_2910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1037_inst_ack_1, ack => convTranspose_CP_814_elements(240)); -- 
    -- CP-element group 241:  join  transition  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	239 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_271/forx_xbody228_forx_xbody228_PhiReq/$exit
      -- CP-element group 241: 	 branch_block_stmt_271/forx_xbody228_forx_xbody228_PhiReq/phi_stmt_1031/$exit
      -- CP-element group 241: 	 branch_block_stmt_271/forx_xbody228_forx_xbody228_PhiReq/phi_stmt_1031/phi_stmt_1031_sources/$exit
      -- CP-element group 241: 	 branch_block_stmt_271/forx_xbody228_forx_xbody228_PhiReq/phi_stmt_1031/phi_stmt_1031_sources/type_cast_1037/$exit
      -- CP-element group 241: 	 branch_block_stmt_271/forx_xbody228_forx_xbody228_PhiReq/phi_stmt_1031/phi_stmt_1031_sources/type_cast_1037/SplitProtocol/$exit
      -- CP-element group 241: 	 branch_block_stmt_271/forx_xbody228_forx_xbody228_PhiReq/phi_stmt_1031/phi_stmt_1031_req
      -- 
    phi_stmt_1031_req_2911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1031_req_2911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(241), ack => phi_stmt_1031_req_1); -- 
    convTranspose_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_814_elements(239) & convTranspose_CP_814_elements(240);
      gj_convTranspose_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_814_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  merge  transition  place  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: 	238 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (2) 
      -- CP-element group 242: 	 branch_block_stmt_271/merge_stmt_1030_PhiReqMerge
      -- CP-element group 242: 	 branch_block_stmt_271/merge_stmt_1030_PhiAck/$entry
      -- 
    convTranspose_CP_814_elements(242) <= OrReduce(convTranspose_CP_814_elements(241) & convTranspose_CP_814_elements(238));
    -- CP-element group 243:  fork  transition  place  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	179 
    -- CP-element group 243: 	180 
    -- CP-element group 243: 	182 
    -- CP-element group 243: 	184 
    -- CP-element group 243:  members (29) 
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061__entry__
      -- CP-element group 243: 	 branch_block_stmt_271/merge_stmt_1030__exit__
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/$entry
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/addr_of_1044_update_start_
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_index_resized_1
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_index_scaled_1
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_index_computed_1
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_index_resize_1/$entry
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_index_resize_1/$exit
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_index_resize_1/index_resize_req
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_index_resize_1/index_resize_ack
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_index_scale_1/$entry
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_index_scale_1/$exit
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_index_scale_1/scale_rename_req
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_index_scale_1/scale_rename_ack
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_final_index_sum_regn_update_start
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_final_index_sum_regn_Sample/$entry
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_final_index_sum_regn_Sample/req
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_final_index_sum_regn_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/array_obj_ref_1043_final_index_sum_regn_Update/req
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/addr_of_1044_complete/$entry
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/addr_of_1044_complete/req
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_update_start_
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_Update/word_access_complete/$entry
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_Update/word_access_complete/word_0/$entry
      -- CP-element group 243: 	 branch_block_stmt_271/assign_stmt_1045_to_assign_stmt_1061/ptr_deref_1047_Update/word_access_complete/word_0/cr
      -- CP-element group 243: 	 branch_block_stmt_271/merge_stmt_1030_PhiAck/$exit
      -- CP-element group 243: 	 branch_block_stmt_271/merge_stmt_1030_PhiAck/phi_stmt_1031_ack
      -- 
    phi_stmt_1031_ack_2916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1031_ack_0, ack => convTranspose_CP_814_elements(243)); -- 
    req_2249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(243), ack => array_obj_ref_1043_index_offset_req_0); -- 
    req_2254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(243), ack => array_obj_ref_1043_index_offset_req_1); -- 
    req_2269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(243), ack => addr_of_1044_final_reg_req_1); -- 
    cr_2319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(243), ack => ptr_deref_1047_store_0_req_1); -- 
    -- CP-element group 244:  merge  fork  transition  place  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	186 
    -- CP-element group 244: 	176 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	188 
    -- CP-element group 244: 	189 
    -- CP-element group 244:  members (13) 
      -- CP-element group 244: 	 branch_block_stmt_271/call_stmt_1072__entry__
      -- CP-element group 244: 	 branch_block_stmt_271/merge_stmt_1070__exit__
      -- CP-element group 244: 	 branch_block_stmt_271/call_stmt_1072/call_stmt_1072_Sample/crr
      -- CP-element group 244: 	 branch_block_stmt_271/call_stmt_1072/call_stmt_1072_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_271/call_stmt_1072/call_stmt_1072_Sample/$entry
      -- CP-element group 244: 	 branch_block_stmt_271/call_stmt_1072/call_stmt_1072_Update/$entry
      -- CP-element group 244: 	 branch_block_stmt_271/call_stmt_1072/call_stmt_1072_update_start_
      -- CP-element group 244: 	 branch_block_stmt_271/call_stmt_1072/call_stmt_1072_Update/ccr
      -- CP-element group 244: 	 branch_block_stmt_271/call_stmt_1072/$entry
      -- CP-element group 244: 	 branch_block_stmt_271/merge_stmt_1070_PhiReqMerge
      -- CP-element group 244: 	 branch_block_stmt_271/merge_stmt_1070_PhiAck/$entry
      -- CP-element group 244: 	 branch_block_stmt_271/merge_stmt_1070_PhiAck/$exit
      -- CP-element group 244: 	 branch_block_stmt_271/merge_stmt_1070_PhiAck/dummy
      -- 
    crr_2350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(244), ack => call_stmt_1072_call_req_0); -- 
    ccr_2355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(244), ack => call_stmt_1072_call_req_1); -- 
    convTranspose_CP_814_elements(244) <= OrReduce(convTranspose_CP_814_elements(186) & convTranspose_CP_814_elements(176));
    -- CP-element group 245:  transition  output  delay-element  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	189 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	248 
    -- CP-element group 245:  members (4) 
      -- CP-element group 245: 	 branch_block_stmt_271/forx_xend235_whilex_xbody_PhiReq/phi_stmt_1098/$exit
      -- CP-element group 245: 	 branch_block_stmt_271/forx_xend235_whilex_xbody_PhiReq/phi_stmt_1098/phi_stmt_1098_sources/$exit
      -- CP-element group 245: 	 branch_block_stmt_271/forx_xend235_whilex_xbody_PhiReq/phi_stmt_1098/phi_stmt_1098_sources/type_cast_1102_konst_delay_trans
      -- CP-element group 245: 	 branch_block_stmt_271/forx_xend235_whilex_xbody_PhiReq/phi_stmt_1098/phi_stmt_1098_req
      -- 
    phi_stmt_1098_req_2950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1098_req_2950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(245), ack => phi_stmt_1098_req_0); -- 
    -- Element group convTranspose_CP_814_elements(245) is a control-delay.
    cp_element_245_delay: control_delay_element  generic map(name => " 245_delay", delay_value => 1)  port map(req => convTranspose_CP_814_elements(189), ack => convTranspose_CP_814_elements(245), clk => clk, reset =>reset);
    -- CP-element group 246:  transition  output  delay-element  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	189 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (4) 
      -- CP-element group 246: 	 branch_block_stmt_271/forx_xend235_whilex_xbody_PhiReq/phi_stmt_1105/$exit
      -- CP-element group 246: 	 branch_block_stmt_271/forx_xend235_whilex_xbody_PhiReq/phi_stmt_1105/phi_stmt_1105_sources/$exit
      -- CP-element group 246: 	 branch_block_stmt_271/forx_xend235_whilex_xbody_PhiReq/phi_stmt_1105/phi_stmt_1105_sources/type_cast_1109_konst_delay_trans
      -- CP-element group 246: 	 branch_block_stmt_271/forx_xend235_whilex_xbody_PhiReq/phi_stmt_1105/phi_stmt_1105_req
      -- 
    phi_stmt_1105_req_2958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1105_req_2958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(246), ack => phi_stmt_1105_req_0); -- 
    -- Element group convTranspose_CP_814_elements(246) is a control-delay.
    cp_element_246_delay: control_delay_element  generic map(name => " 246_delay", delay_value => 1)  port map(req => convTranspose_CP_814_elements(189), ack => convTranspose_CP_814_elements(246), clk => clk, reset =>reset);
    -- CP-element group 247:  transition  output  delay-element  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	189 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (4) 
      -- CP-element group 247: 	 branch_block_stmt_271/forx_xend235_whilex_xbody_PhiReq/phi_stmt_1112/$exit
      -- CP-element group 247: 	 branch_block_stmt_271/forx_xend235_whilex_xbody_PhiReq/phi_stmt_1112/phi_stmt_1112_sources/$exit
      -- CP-element group 247: 	 branch_block_stmt_271/forx_xend235_whilex_xbody_PhiReq/phi_stmt_1112/phi_stmt_1112_sources/type_cast_1116_konst_delay_trans
      -- CP-element group 247: 	 branch_block_stmt_271/forx_xend235_whilex_xbody_PhiReq/phi_stmt_1112/phi_stmt_1112_req
      -- 
    phi_stmt_1112_req_2966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1112_req_2966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(247), ack => phi_stmt_1112_req_0); -- 
    -- Element group convTranspose_CP_814_elements(247) is a control-delay.
    cp_element_247_delay: control_delay_element  generic map(name => " 247_delay", delay_value => 1)  port map(req => convTranspose_CP_814_elements(189), ack => convTranspose_CP_814_elements(247), clk => clk, reset =>reset);
    -- CP-element group 248:  join  transition  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: 	245 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	259 
    -- CP-element group 248:  members (1) 
      -- CP-element group 248: 	 branch_block_stmt_271/forx_xend235_whilex_xbody_PhiReq/$exit
      -- 
    convTranspose_cp_element_group_248: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_248"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_814_elements(247) & convTranspose_CP_814_elements(245) & convTranspose_CP_814_elements(246);
      gj_convTranspose_cp_element_group_248 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_814_elements(248), clk => clk, reset => reset); --
    end block;
    -- CP-element group 249:  transition  input  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	213 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	251 
    -- CP-element group 249:  members (2) 
      -- CP-element group 249: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1098/phi_stmt_1098_sources/type_cast_1104/SplitProtocol/Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1098/phi_stmt_1098_sources/type_cast_1104/SplitProtocol/Sample/ra
      -- 
    ra_2986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1104_inst_ack_0, ack => convTranspose_CP_814_elements(249)); -- 
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	213 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (2) 
      -- CP-element group 250: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1098/phi_stmt_1098_sources/type_cast_1104/SplitProtocol/Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1098/phi_stmt_1098_sources/type_cast_1104/SplitProtocol/Update/ca
      -- 
    ca_2991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1104_inst_ack_1, ack => convTranspose_CP_814_elements(250)); -- 
    -- CP-element group 251:  join  transition  output  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	258 
    -- CP-element group 251:  members (5) 
      -- CP-element group 251: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1098/$exit
      -- CP-element group 251: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1098/phi_stmt_1098_sources/$exit
      -- CP-element group 251: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1098/phi_stmt_1098_sources/type_cast_1104/$exit
      -- CP-element group 251: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1098/phi_stmt_1098_sources/type_cast_1104/SplitProtocol/$exit
      -- CP-element group 251: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1098/phi_stmt_1098_req
      -- 
    phi_stmt_1098_req_2992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1098_req_2992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(251), ack => phi_stmt_1098_req_1); -- 
    convTranspose_cp_element_group_251: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_251"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_814_elements(249) & convTranspose_CP_814_elements(250);
      gj_convTranspose_cp_element_group_251 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_814_elements(251), clk => clk, reset => reset); --
    end block;
    -- CP-element group 252:  transition  input  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	213 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	254 
    -- CP-element group 252:  members (2) 
      -- CP-element group 252: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1105/phi_stmt_1105_sources/type_cast_1111/SplitProtocol/Sample/$exit
      -- CP-element group 252: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1105/phi_stmt_1105_sources/type_cast_1111/SplitProtocol/Sample/ra
      -- 
    ra_3009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1111_inst_ack_0, ack => convTranspose_CP_814_elements(252)); -- 
    -- CP-element group 253:  transition  input  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	213 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (2) 
      -- CP-element group 253: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1105/phi_stmt_1105_sources/type_cast_1111/SplitProtocol/Update/$exit
      -- CP-element group 253: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1105/phi_stmt_1105_sources/type_cast_1111/SplitProtocol/Update/ca
      -- 
    ca_3014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1111_inst_ack_1, ack => convTranspose_CP_814_elements(253)); -- 
    -- CP-element group 254:  join  transition  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	252 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	258 
    -- CP-element group 254:  members (5) 
      -- CP-element group 254: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1105/$exit
      -- CP-element group 254: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1105/phi_stmt_1105_sources/$exit
      -- CP-element group 254: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1105/phi_stmt_1105_sources/type_cast_1111/$exit
      -- CP-element group 254: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1105/phi_stmt_1105_sources/type_cast_1111/SplitProtocol/$exit
      -- CP-element group 254: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1105/phi_stmt_1105_req
      -- 
    phi_stmt_1105_req_3015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1105_req_3015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(254), ack => phi_stmt_1105_req_1); -- 
    convTranspose_cp_element_group_254: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_254"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_814_elements(252) & convTranspose_CP_814_elements(253);
      gj_convTranspose_cp_element_group_254 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_814_elements(254), clk => clk, reset => reset); --
    end block;
    -- CP-element group 255:  transition  input  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	213 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	257 
    -- CP-element group 255:  members (2) 
      -- CP-element group 255: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1112/phi_stmt_1112_sources/type_cast_1118/SplitProtocol/Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1112/phi_stmt_1112_sources/type_cast_1118/SplitProtocol/Sample/ra
      -- 
    ra_3032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1118_inst_ack_0, ack => convTranspose_CP_814_elements(255)); -- 
    -- CP-element group 256:  transition  input  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	213 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (2) 
      -- CP-element group 256: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1112/phi_stmt_1112_sources/type_cast_1118/SplitProtocol/Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1112/phi_stmt_1112_sources/type_cast_1118/SplitProtocol/Update/ca
      -- 
    ca_3037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1118_inst_ack_1, ack => convTranspose_CP_814_elements(256)); -- 
    -- CP-element group 257:  join  transition  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: 	255 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (5) 
      -- CP-element group 257: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1112/$exit
      -- CP-element group 257: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1112/phi_stmt_1112_sources/$exit
      -- CP-element group 257: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1112/phi_stmt_1112_sources/type_cast_1118/$exit
      -- CP-element group 257: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1112/phi_stmt_1112_sources/type_cast_1118/SplitProtocol/$exit
      -- CP-element group 257: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1112/phi_stmt_1112_req
      -- 
    phi_stmt_1112_req_3038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1112_req_3038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(257), ack => phi_stmt_1112_req_1); -- 
    convTranspose_cp_element_group_257: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_257"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_814_elements(256) & convTranspose_CP_814_elements(255);
      gj_convTranspose_cp_element_group_257 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_814_elements(257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 258:  join  transition  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	251 
    -- CP-element group 258: 	257 
    -- CP-element group 258: 	254 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (1) 
      -- CP-element group 258: 	 branch_block_stmt_271/whilex_xbody_whilex_xbody_PhiReq/$exit
      -- 
    convTranspose_cp_element_group_258: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_258"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_814_elements(251) & convTranspose_CP_814_elements(257) & convTranspose_CP_814_elements(254);
      gj_convTranspose_cp_element_group_258 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_814_elements(258), clk => clk, reset => reset); --
    end block;
    -- CP-element group 259:  merge  fork  transition  place  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	248 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259: 	261 
    -- CP-element group 259: 	262 
    -- CP-element group 259:  members (2) 
      -- CP-element group 259: 	 branch_block_stmt_271/merge_stmt_1097_PhiReqMerge
      -- CP-element group 259: 	 branch_block_stmt_271/merge_stmt_1097_PhiAck/$entry
      -- 
    convTranspose_CP_814_elements(259) <= OrReduce(convTranspose_CP_814_elements(248) & convTranspose_CP_814_elements(258));
    -- CP-element group 260:  transition  input  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	263 
    -- CP-element group 260:  members (1) 
      -- CP-element group 260: 	 branch_block_stmt_271/merge_stmt_1097_PhiAck/phi_stmt_1098_ack
      -- 
    phi_stmt_1098_ack_3043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1098_ack_0, ack => convTranspose_CP_814_elements(260)); -- 
    -- CP-element group 261:  transition  input  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	259 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	263 
    -- CP-element group 261:  members (1) 
      -- CP-element group 261: 	 branch_block_stmt_271/merge_stmt_1097_PhiAck/phi_stmt_1105_ack
      -- 
    phi_stmt_1105_ack_3044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1105_ack_0, ack => convTranspose_CP_814_elements(261)); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	259 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	263 
    -- CP-element group 262:  members (1) 
      -- CP-element group 262: 	 branch_block_stmt_271/merge_stmt_1097_PhiAck/phi_stmt_1112_ack
      -- 
    phi_stmt_1112_ack_3045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1112_ack_0, ack => convTranspose_CP_814_elements(262)); -- 
    -- CP-element group 263:  join  fork  transition  place  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	260 
    -- CP-element group 263: 	261 
    -- CP-element group 263: 	262 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	190 
    -- CP-element group 263: 	206 
    -- CP-element group 263: 	207 
    -- CP-element group 263: 	208 
    -- CP-element group 263: 	191 
    -- CP-element group 263: 	197 
    -- CP-element group 263: 	201 
    -- CP-element group 263: 	203 
    -- CP-element group 263: 	193 
    -- CP-element group 263: 	195 
    -- CP-element group 263: 	198 
    -- CP-element group 263: 	199 
    -- CP-element group 263: 	210 
    -- CP-element group 263:  members (47) 
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274__entry__
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_Update/word_access_complete/$entry
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_Update/word_access_complete/word_0/$entry
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1195_complete/$entry
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1235_update_start_
      -- CP-element group 263: 	 branch_block_stmt_271/merge_stmt_1097__exit__
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_Update/word_access_complete/word_0/cr
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1235_Update/cr
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1235_sample_start_
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_final_index_sum_regn_Update/req
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_update_start_
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1195_complete/req
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_Update/word_access_complete/word_0/$entry
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_final_index_sum_regn_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1235_Sample/$entry
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1216_complete/$entry
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1216_complete/req
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1235_Sample/rr
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_update_start_
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_Update/word_access_complete/$entry
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1235_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1215_final_index_sum_regn_update_start
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_final_index_sum_regn_Update/req
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_final_index_sum_regn_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1219_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1216_update_start_
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/addr_of_1195_update_start_
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1203_Update/cr
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1182_Update/cr
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1182_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1256_Update/cr
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1256_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/$entry
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1203_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1182_Sample/rr
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1182_Sample/$entry
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1182_update_start_
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1182_sample_start_
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1203_Sample/rr
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1203_Sample/$entry
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/array_obj_ref_1194_final_index_sum_regn_update_start
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1203_update_start_
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1256_update_start_
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/type_cast_1203_sample_start_
      -- CP-element group 263: 	 branch_block_stmt_271/assign_stmt_1124_to_assign_stmt_1274/ptr_deref_1199_Update/word_access_complete/word_0/cr
      -- CP-element group 263: 	 branch_block_stmt_271/merge_stmt_1097_PhiAck/$exit
      -- 
    cr_2581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(263), ack => ptr_deref_1219_store_0_req_1); -- 
    cr_2595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(263), ack => type_cast_1235_inst_req_1); -- 
    req_2516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(263), ack => array_obj_ref_1215_index_offset_req_1); -- 
    req_2421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(263), ack => addr_of_1195_final_reg_req_1); -- 
    req_2531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(263), ack => addr_of_1216_final_reg_req_1); -- 
    rr_2590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(263), ack => type_cast_1235_inst_req_0); -- 
    req_2406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(263), ack => array_obj_ref_1194_index_offset_req_1); -- 
    cr_2485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(263), ack => type_cast_1203_inst_req_1); -- 
    cr_2375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(263), ack => type_cast_1182_inst_req_1); -- 
    cr_2609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(263), ack => type_cast_1256_inst_req_1); -- 
    rr_2370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(263), ack => type_cast_1182_inst_req_0); -- 
    rr_2480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(263), ack => type_cast_1203_inst_req_0); -- 
    cr_2466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_814_elements(263), ack => ptr_deref_1199_load_0_req_1); -- 
    convTranspose_cp_element_group_263: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_263"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_814_elements(260) & convTranspose_CP_814_elements(261) & convTranspose_CP_814_elements(262);
      gj_convTranspose_cp_element_group_263 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_814_elements(263), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar402_723_resized : std_logic_vector(13 downto 0);
    signal R_indvar402_723_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1042_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1042_scaled : std_logic_vector(13 downto 0);
    signal R_shr307364_1193_resized : std_logic_vector(13 downto 0);
    signal R_shr307364_1193_scaled : std_logic_vector(13 downto 0);
    signal R_shr313366_1214_resized : std_logic_vector(13 downto 0);
    signal R_shr313366_1214_scaled : std_logic_vector(13 downto 0);
    signal add105_547 : std_logic_vector(15 downto 0);
    signal add114_572 : std_logic_vector(15 downto 0);
    signal add123_597 : std_logic_vector(15 downto 0);
    signal add13_322 : std_logic_vector(31 downto 0);
    signal add167_751 : std_logic_vector(63 downto 0);
    signal add173_769 : std_logic_vector(63 downto 0);
    signal add179_787 : std_logic_vector(63 downto 0);
    signal add185_805 : std_logic_vector(63 downto 0);
    signal add191_823 : std_logic_vector(63 downto 0);
    signal add197_841 : std_logic_vector(63 downto 0);
    signal add203_859 : std_logic_vector(63 downto 0);
    signal add23_347 : std_logic_vector(15 downto 0);
    signal add257_1079 : std_logic_vector(15 downto 0);
    signal add269_1090 : std_logic_vector(15 downto 0);
    signal add286_1144 : std_logic_vector(15 downto 0);
    signal add288_1154 : std_logic_vector(15 downto 0);
    signal add301_1169 : std_logic_vector(15 downto 0);
    signal add303_1179 : std_logic_vector(15 downto 0);
    signal add318_1227 : std_logic_vector(15 downto 0);
    signal add33_372 : std_logic_vector(15 downto 0);
    signal add43_397 : std_logic_vector(15 downto 0);
    signal add53_422 : std_logic_vector(15 downto 0);
    signal add66_447 : std_logic_vector(31 downto 0);
    signal add75_472 : std_logic_vector(15 downto 0);
    signal add84_497 : std_logic_vector(15 downto 0);
    signal add93_522 : std_logic_vector(31 downto 0);
    signal add_297 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1043_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1043_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1043_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1043_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1043_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1043_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1194_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1194_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1194_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1194_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1194_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1194_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1215_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1215_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1215_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1215_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1215_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1215_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_724_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_724_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_724_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_724_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_724_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_724_root_address : std_logic_vector(13 downto 0);
    signal arrayidx231_1045 : std_logic_vector(31 downto 0);
    signal arrayidx309_1196 : std_logic_vector(31 downto 0);
    signal arrayidx315_1217 : std_logic_vector(31 downto 0);
    signal arrayidx_726 : std_logic_vector(31 downto 0);
    signal call103_538 : std_logic_vector(7 downto 0);
    signal call107_550 : std_logic_vector(7 downto 0);
    signal call112_563 : std_logic_vector(7 downto 0);
    signal call116_575 : std_logic_vector(7 downto 0);
    signal call11_313 : std_logic_vector(7 downto 0);
    signal call121_588 : std_logic_vector(7 downto 0);
    signal call160_729 : std_logic_vector(7 downto 0);
    signal call164_742 : std_logic_vector(7 downto 0);
    signal call16_325 : std_logic_vector(7 downto 0);
    signal call170_760 : std_logic_vector(7 downto 0);
    signal call176_778 : std_logic_vector(7 downto 0);
    signal call182_796 : std_logic_vector(7 downto 0);
    signal call188_814 : std_logic_vector(7 downto 0);
    signal call194_832 : std_logic_vector(7 downto 0);
    signal call200_850 : std_logic_vector(7 downto 0);
    signal call21_338 : std_logic_vector(7 downto 0);
    signal call237_1072 : std_logic_vector(63 downto 0);
    signal call26_350 : std_logic_vector(7 downto 0);
    signal call2_288 : std_logic_vector(7 downto 0);
    signal call31_363 : std_logic_vector(7 downto 0);
    signal call348_1290 : std_logic_vector(63 downto 0);
    signal call36_375 : std_logic_vector(7 downto 0);
    signal call41_388 : std_logic_vector(7 downto 0);
    signal call46_400 : std_logic_vector(7 downto 0);
    signal call51_413 : std_logic_vector(7 downto 0);
    signal call59_425 : std_logic_vector(7 downto 0);
    signal call64_438 : std_logic_vector(7 downto 0);
    signal call68_450 : std_logic_vector(7 downto 0);
    signal call6_300 : std_logic_vector(7 downto 0);
    signal call73_463 : std_logic_vector(7 downto 0);
    signal call77_475 : std_logic_vector(7 downto 0);
    signal call82_488 : std_logic_vector(7 downto 0);
    signal call86_500 : std_logic_vector(7 downto 0);
    signal call91_513 : std_logic_vector(7 downto 0);
    signal call98_525 : std_logic_vector(7 downto 0);
    signal call_274 : std_logic_vector(7 downto 0);
    signal cmp212372_890 : std_logic_vector(0 downto 0);
    signal cmp226369_986 : std_logic_vector(0 downto 0);
    signal cmp324_1232 : std_logic_vector(0 downto 0);
    signal cmp332_1253 : std_logic_vector(0 downto 0);
    signal cmp342_1274 : std_logic_vector(0 downto 0);
    signal cmp376_667 : std_logic_vector(0 downto 0);
    signal conv101_529 : std_logic_vector(15 downto 0);
    signal conv104_542 : std_logic_vector(15 downto 0);
    signal conv110_554 : std_logic_vector(15 downto 0);
    signal conv113_567 : std_logic_vector(15 downto 0);
    signal conv119_579 : std_logic_vector(15 downto 0);
    signal conv122_592 : std_logic_vector(15 downto 0);
    signal conv128_602 : std_logic_vector(31 downto 0);
    signal conv12_317 : std_logic_vector(31 downto 0);
    signal conv130_606 : std_logic_vector(31 downto 0);
    signal conv132_610 : std_logic_vector(31 downto 0);
    signal conv138_624 : std_logic_vector(31 downto 0);
    signal conv141_628 : std_logic_vector(31 downto 0);
    signal conv147_642 : std_logic_vector(31 downto 0);
    signal conv150_646 : std_logic_vector(31 downto 0);
    signal conv161_733 : std_logic_vector(63 downto 0);
    signal conv166_746 : std_logic_vector(63 downto 0);
    signal conv172_764 : std_logic_vector(63 downto 0);
    signal conv178_782 : std_logic_vector(63 downto 0);
    signal conv184_800 : std_logic_vector(63 downto 0);
    signal conv190_818 : std_logic_vector(63 downto 0);
    signal conv196_836 : std_logic_vector(63 downto 0);
    signal conv19_329 : std_logic_vector(15 downto 0);
    signal conv1_279 : std_logic_vector(15 downto 0);
    signal conv202_854 : std_logic_vector(63 downto 0);
    signal conv22_342 : std_logic_vector(15 downto 0);
    signal conv238_1287 : std_logic_vector(63 downto 0);
    signal conv29_354 : std_logic_vector(15 downto 0);
    signal conv306_1183 : std_logic_vector(63 downto 0);
    signal conv312_1204 : std_logic_vector(63 downto 0);
    signal conv32_367 : std_logic_vector(15 downto 0);
    signal conv349_1295 : std_logic_vector(63 downto 0);
    signal conv39_379 : std_logic_vector(15 downto 0);
    signal conv3_292 : std_logic_vector(15 downto 0);
    signal conv42_392 : std_logic_vector(15 downto 0);
    signal conv49_404 : std_logic_vector(15 downto 0);
    signal conv52_417 : std_logic_vector(15 downto 0);
    signal conv62_429 : std_logic_vector(31 downto 0);
    signal conv65_442 : std_logic_vector(31 downto 0);
    signal conv71_454 : std_logic_vector(15 downto 0);
    signal conv74_467 : std_logic_vector(15 downto 0);
    signal conv80_479 : std_logic_vector(15 downto 0);
    signal conv83_492 : std_logic_vector(15 downto 0);
    signal conv89_504 : std_logic_vector(31 downto 0);
    signal conv92_517 : std_logic_vector(31 downto 0);
    signal conv9_304 : std_logic_vector(31 downto 0);
    signal exitcond1_1061 : std_logic_vector(0 downto 0);
    signal exitcond2_874 : std_logic_vector(0 downto 0);
    signal exitcond_970 : std_logic_vector(0 downto 0);
    signal iNsTr_27_696 : std_logic_vector(63 downto 0);
    signal iNsTr_40_934 : std_logic_vector(63 downto 0);
    signal iNsTr_44_950 : std_logic_vector(63 downto 0);
    signal iNsTr_47_1015 : std_logic_vector(63 downto 0);
    signal inc327_1236 : std_logic_vector(15 downto 0);
    signal inc327x_xinput_dim1x_x1_1241 : std_logic_vector(15 downto 0);
    signal inc336_1257 : std_logic_vector(15 downto 0);
    signal inc336x_xinput_dim0x_x1_1262 : std_logic_vector(15 downto 0);
    signal indvar402_712 : std_logic_vector(63 downto 0);
    signal indvar_1031 : std_logic_vector(63 downto 0);
    signal indvarx_xnext389_965 : std_logic_vector(63 downto 0);
    signal indvarx_xnext403_869 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1056 : std_logic_vector(63 downto 0);
    signal input_dim0x_x1_1098 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1105 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1269 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0_1112 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1248 : std_logic_vector(15 downto 0);
    signal mul133_620 : std_logic_vector(31 downto 0);
    signal mul139_633 : std_logic_vector(31 downto 0);
    signal mul142_638 : std_logic_vector(31 downto 0);
    signal mul148_651 : std_logic_vector(31 downto 0);
    signal mul151_656 : std_logic_vector(31 downto 0);
    signal mul154_661 : std_logic_vector(31 downto 0);
    signal mul254_1124 : std_logic_vector(15 downto 0);
    signal mul266_1134 : std_logic_vector(15 downto 0);
    signal mul285_1139 : std_logic_vector(15 downto 0);
    signal mul287_1149 : std_logic_vector(15 downto 0);
    signal mul300_1159 : std_logic_vector(15 downto 0);
    signal mul302_1174 : std_logic_vector(15 downto 0);
    signal mul_615 : std_logic_vector(31 downto 0);
    signal ptr_deref_1047_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1047_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1047_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1047_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1047_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1047_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1199_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1199_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1199_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1199_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1199_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1219_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1219_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1219_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1219_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1219_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1219_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_861_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_861_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_861_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_861_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_861_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_861_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl102_535 : std_logic_vector(15 downto 0);
    signal shl10_310 : std_logic_vector(31 downto 0);
    signal shl111_560 : std_logic_vector(15 downto 0);
    signal shl120_585 : std_logic_vector(15 downto 0);
    signal shl163_739 : std_logic_vector(63 downto 0);
    signal shl169_757 : std_logic_vector(63 downto 0);
    signal shl175_775 : std_logic_vector(63 downto 0);
    signal shl181_793 : std_logic_vector(63 downto 0);
    signal shl187_811 : std_logic_vector(63 downto 0);
    signal shl193_829 : std_logic_vector(63 downto 0);
    signal shl199_847 : std_logic_vector(63 downto 0);
    signal shl20_335 : std_logic_vector(15 downto 0);
    signal shl30_360 : std_logic_vector(15 downto 0);
    signal shl40_385 : std_logic_vector(15 downto 0);
    signal shl50_410 : std_logic_vector(15 downto 0);
    signal shl63_435 : std_logic_vector(31 downto 0);
    signal shl72_460 : std_logic_vector(15 downto 0);
    signal shl81_485 : std_logic_vector(15 downto 0);
    signal shl90_510 : std_logic_vector(31 downto 0);
    signal shl_285 : std_logic_vector(15 downto 0);
    signal shr307364_1189 : std_logic_vector(63 downto 0);
    signal shr313366_1210 : std_logic_vector(63 downto 0);
    signal sub260_1129 : std_logic_vector(15 downto 0);
    signal sub272_1095 : std_logic_vector(15 downto 0);
    signal sub273_1164 : std_logic_vector(15 downto 0);
    signal sub353_1300 : std_logic_vector(63 downto 0);
    signal sub_1084 : std_logic_vector(15 downto 0);
    signal tmp310_1200 : std_logic_vector(63 downto 0);
    signal tmp383_999 : std_logic_vector(31 downto 0);
    signal tmp383x_xop_1011 : std_logic_vector(31 downto 0);
    signal tmp384_1005 : std_logic_vector(0 downto 0);
    signal tmp387_1028 : std_logic_vector(63 downto 0);
    signal tmp390_902 : std_logic_vector(31 downto 0);
    signal tmp392_907 : std_logic_vector(31 downto 0);
    signal tmp394_912 : std_logic_vector(31 downto 0);
    signal tmp395_918 : std_logic_vector(31 downto 0);
    signal tmp395x_xop_930 : std_logic_vector(31 downto 0);
    signal tmp396_924 : std_logic_vector(0 downto 0);
    signal tmp400_947 : std_logic_vector(63 downto 0);
    signal tmp409_680 : std_logic_vector(31 downto 0);
    signal tmp409x_xop_692 : std_logic_vector(31 downto 0);
    signal tmp410_686 : std_logic_vector(0 downto 0);
    signal tmp414_709 : std_logic_vector(63 downto 0);
    signal type_cast_1003_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1009_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1019_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1026_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1035_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1037_wire : std_logic_vector(63 downto 0);
    signal type_cast_1049_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1054_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1077_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1088_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1102_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1104_wire : std_logic_vector(15 downto 0);
    signal type_cast_1109_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1111_wire : std_logic_vector(15 downto 0);
    signal type_cast_1116_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1118_wire : std_logic_vector(15 downto 0);
    signal type_cast_1187_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1208_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1225_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1245_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1266_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1285_wire : std_logic_vector(63 downto 0);
    signal type_cast_1293_wire : std_logic_vector(63 downto 0);
    signal type_cast_283_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_308_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_333_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_358_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_383_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_408_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_433_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_458_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_483_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_508_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_533_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_558_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_583_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_665_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_678_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_684_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_690_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_700_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_707_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_716_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_718_wire : std_logic_vector(63 downto 0);
    signal type_cast_737_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_755_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_773_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_791_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_809_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_827_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_845_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_867_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_888_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_916_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_922_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_928_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_938_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_945_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_954_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_956_wire : std_logic_vector(63 downto 0);
    signal type_cast_963_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_984_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_997_wire_constant : std_logic_vector(31 downto 0);
    signal xx_xop416_940 : std_logic_vector(63 downto 0);
    signal xx_xop417_702 : std_logic_vector(63 downto 0);
    signal xx_xop_1021 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1043_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1043_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1043_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1043_resized_base_address <= "00000000000000";
    array_obj_ref_1194_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1194_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1194_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1194_resized_base_address <= "00000000000000";
    array_obj_ref_1215_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1215_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1215_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1215_resized_base_address <= "00000000000000";
    array_obj_ref_724_constant_part_of_offset <= "00000000000000";
    array_obj_ref_724_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_724_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_724_resized_base_address <= "00000000000000";
    ptr_deref_1047_word_offset_0 <= "00000000000000";
    ptr_deref_1199_word_offset_0 <= "00000000000000";
    ptr_deref_1219_word_offset_0 <= "00000000000000";
    ptr_deref_861_word_offset_0 <= "00000000000000";
    type_cast_1003_wire_constant <= "00000000000000000000000000000001";
    type_cast_1009_wire_constant <= "11111111111111111111111111111111";
    type_cast_1019_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1026_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1035_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1049_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1054_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1077_wire_constant <= "1111111111111111";
    type_cast_1088_wire_constant <= "1111111111111111";
    type_cast_1102_wire_constant <= "0000000000000000";
    type_cast_1109_wire_constant <= "0000000000000000";
    type_cast_1116_wire_constant <= "0000000000000000";
    type_cast_1187_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1208_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1225_wire_constant <= "0000000000000100";
    type_cast_1245_wire_constant <= "0000000000000000";
    type_cast_1266_wire_constant <= "0000000000000000";
    type_cast_283_wire_constant <= "0000000000001000";
    type_cast_308_wire_constant <= "00000000000000000000000000001000";
    type_cast_333_wire_constant <= "0000000000001000";
    type_cast_358_wire_constant <= "0000000000001000";
    type_cast_383_wire_constant <= "0000000000001000";
    type_cast_408_wire_constant <= "0000000000001000";
    type_cast_433_wire_constant <= "00000000000000000000000000001000";
    type_cast_458_wire_constant <= "0000000000001000";
    type_cast_483_wire_constant <= "0000000000001000";
    type_cast_508_wire_constant <= "00000000000000000000000000001000";
    type_cast_533_wire_constant <= "0000000000001000";
    type_cast_558_wire_constant <= "0000000000001000";
    type_cast_583_wire_constant <= "0000000000001000";
    type_cast_665_wire_constant <= "00000000000000000000000000000011";
    type_cast_678_wire_constant <= "00000000000000000000000000000010";
    type_cast_684_wire_constant <= "00000000000000000000000000000001";
    type_cast_690_wire_constant <= "11111111111111111111111111111111";
    type_cast_700_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_707_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_716_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_737_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_755_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_773_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_791_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_809_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_827_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_845_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_867_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_888_wire_constant <= "00000000000000000000000000000011";
    type_cast_916_wire_constant <= "00000000000000000000000000000010";
    type_cast_922_wire_constant <= "00000000000000000000000000000001";
    type_cast_928_wire_constant <= "11111111111111111111111111111111";
    type_cast_938_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_945_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_954_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_963_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_984_wire_constant <= "00000000000000000000000000000011";
    type_cast_997_wire_constant <= "00000000000000000000000000000010";
    phi_stmt_1031: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1035_wire_constant & type_cast_1037_wire;
      req <= phi_stmt_1031_req_0 & phi_stmt_1031_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1031",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1031_ack_0,
          idata => idata,
          odata => indvar_1031,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1031
    phi_stmt_1098: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1102_wire_constant & type_cast_1104_wire;
      req <= phi_stmt_1098_req_0 & phi_stmt_1098_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1098",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1098_ack_0,
          idata => idata,
          odata => input_dim0x_x1_1098,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1098
    phi_stmt_1105: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1109_wire_constant & type_cast_1111_wire;
      req <= phi_stmt_1105_req_0 & phi_stmt_1105_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1105",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1105_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1105,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1105
    phi_stmt_1112: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1116_wire_constant & type_cast_1118_wire;
      req <= phi_stmt_1112_req_0 & phi_stmt_1112_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1112",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1112_ack_0,
          idata => idata,
          odata => input_dim2x_x0_1112,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1112
    phi_stmt_712: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_716_wire_constant & type_cast_718_wire;
      req <= phi_stmt_712_req_0 & phi_stmt_712_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_712",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_712_ack_0,
          idata => idata,
          odata => indvar402_712,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_712
    phi_stmt_950: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_954_wire_constant & type_cast_956_wire;
      req <= phi_stmt_950_req_0 & phi_stmt_950_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_950",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_950_ack_0,
          idata => idata,
          odata => iNsTr_44_950,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_950
    -- flow-through select operator MUX_1027_inst
    tmp387_1028 <= xx_xop_1021 when (tmp384_1005(0) /=  '0') else type_cast_1026_wire_constant;
    -- flow-through select operator MUX_1247_inst
    input_dim2x_x1_1248 <= type_cast_1245_wire_constant when (cmp324_1232(0) /=  '0') else add318_1227;
    -- flow-through select operator MUX_1268_inst
    input_dim1x_x2_1269 <= type_cast_1266_wire_constant when (cmp332_1253(0) /=  '0') else inc327x_xinput_dim1x_x1_1241;
    -- flow-through select operator MUX_708_inst
    tmp414_709 <= xx_xop417_702 when (tmp410_686(0) /=  '0') else type_cast_707_wire_constant;
    -- flow-through select operator MUX_946_inst
    tmp400_947 <= xx_xop416_940 when (tmp396_924(0) /=  '0') else type_cast_945_wire_constant;
    addr_of_1044_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1044_final_reg_req_0;
      addr_of_1044_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1044_final_reg_req_1;
      addr_of_1044_final_reg_ack_1<= rack(0);
      addr_of_1044_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1044_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1043_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx231_1045,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1195_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1195_final_reg_req_0;
      addr_of_1195_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1195_final_reg_req_1;
      addr_of_1195_final_reg_ack_1<= rack(0);
      addr_of_1195_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1195_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1194_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx309_1196,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1216_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1216_final_reg_req_0;
      addr_of_1216_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1216_final_reg_req_1;
      addr_of_1216_final_reg_ack_1<= rack(0);
      addr_of_1216_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1216_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1215_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx315_1217,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_725_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_725_final_reg_req_0;
      addr_of_725_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_725_final_reg_req_1;
      addr_of_725_final_reg_ack_1<= rack(0);
      addr_of_725_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_725_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_724_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_726,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1014_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1014_inst_req_0;
      type_cast_1014_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1014_inst_req_1;
      type_cast_1014_inst_ack_1<= rack(0);
      type_cast_1014_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1014_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp383x_xop_1011,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_47_1015,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1037_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1037_inst_req_0;
      type_cast_1037_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1037_inst_req_1;
      type_cast_1037_inst_ack_1<= rack(0);
      type_cast_1037_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1037_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1056,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1037_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1104_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1104_inst_req_0;
      type_cast_1104_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1104_inst_req_1;
      type_cast_1104_inst_ack_1<= rack(0);
      type_cast_1104_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1104_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc336x_xinput_dim0x_x1_1262,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1104_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1111_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1111_inst_req_0;
      type_cast_1111_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1111_inst_req_1;
      type_cast_1111_inst_ack_1<= rack(0);
      type_cast_1111_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1111_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1269,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1111_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1118_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1118_inst_req_0;
      type_cast_1118_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1118_inst_req_1;
      type_cast_1118_inst_ack_1<= rack(0);
      type_cast_1118_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1118_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1248,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1118_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1182_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1182_inst_req_0;
      type_cast_1182_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1182_inst_req_1;
      type_cast_1182_inst_ack_1<= rack(0);
      type_cast_1182_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1182_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add288_1154,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv306_1183,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1203_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1203_inst_req_0;
      type_cast_1203_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1203_inst_req_1;
      type_cast_1203_inst_ack_1<= rack(0);
      type_cast_1203_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1203_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add303_1179,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv312_1204,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1235_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1235_inst_req_0;
      type_cast_1235_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1235_inst_req_1;
      type_cast_1235_inst_ack_1<= rack(0);
      type_cast_1235_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1235_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp324_1232,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc327_1236,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1256_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1256_inst_req_0;
      type_cast_1256_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1256_inst_req_1;
      type_cast_1256_inst_ack_1<= rack(0);
      type_cast_1256_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1256_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp332_1253,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc336_1257,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1286_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1286_inst_req_0;
      type_cast_1286_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1286_inst_req_1;
      type_cast_1286_inst_ack_1<= rack(0);
      type_cast_1286_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1286_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1285_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv238_1287,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1294_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1294_inst_req_0;
      type_cast_1294_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1294_inst_req_1;
      type_cast_1294_inst_ack_1<= rack(0);
      type_cast_1294_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1294_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1293_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv349_1295,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_278_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_278_inst_req_0;
      type_cast_278_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_278_inst_req_1;
      type_cast_278_inst_ack_1<= rack(0);
      type_cast_278_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_278_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_274,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_279,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_291_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_291_inst_req_0;
      type_cast_291_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_291_inst_req_1;
      type_cast_291_inst_ack_1<= rack(0);
      type_cast_291_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_291_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_288,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_292,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_303_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_303_inst_req_0;
      type_cast_303_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_303_inst_req_1;
      type_cast_303_inst_ack_1<= rack(0);
      type_cast_303_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_303_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_300,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9_304,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_316_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_316_inst_req_0;
      type_cast_316_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_316_inst_req_1;
      type_cast_316_inst_ack_1<= rack(0);
      type_cast_316_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_316_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call11_313,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_317,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_328_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_328_inst_req_0;
      type_cast_328_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_328_inst_req_1;
      type_cast_328_inst_ack_1<= rack(0);
      type_cast_328_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_328_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_325,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_329,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_341_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_341_inst_req_0;
      type_cast_341_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_341_inst_req_1;
      type_cast_341_inst_ack_1<= rack(0);
      type_cast_341_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_341_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call21_338,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_342,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_353_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_353_inst_req_0;
      type_cast_353_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_353_inst_req_1;
      type_cast_353_inst_ack_1<= rack(0);
      type_cast_353_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_353_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call26_350,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_354,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_366_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_366_inst_req_0;
      type_cast_366_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_366_inst_req_1;
      type_cast_366_inst_ack_1<= rack(0);
      type_cast_366_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_366_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call31_363,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_367,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_378_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_378_inst_req_0;
      type_cast_378_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_378_inst_req_1;
      type_cast_378_inst_ack_1<= rack(0);
      type_cast_378_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_378_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call36_375,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_379,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_391_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_391_inst_req_0;
      type_cast_391_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_391_inst_req_1;
      type_cast_391_inst_ack_1<= rack(0);
      type_cast_391_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_391_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_388,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_392,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_403_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_403_inst_req_0;
      type_cast_403_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_403_inst_req_1;
      type_cast_403_inst_ack_1<= rack(0);
      type_cast_403_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_403_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_400,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv49_404,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_416_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_416_inst_req_0;
      type_cast_416_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_416_inst_req_1;
      type_cast_416_inst_ack_1<= rack(0);
      type_cast_416_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_416_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call51_413,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_417,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_428_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_428_inst_req_0;
      type_cast_428_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_428_inst_req_1;
      type_cast_428_inst_ack_1<= rack(0);
      type_cast_428_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_428_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call59_425,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_429,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_441_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_441_inst_req_0;
      type_cast_441_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_441_inst_req_1;
      type_cast_441_inst_ack_1<= rack(0);
      type_cast_441_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_441_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call64_438,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_442,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_453_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_453_inst_req_0;
      type_cast_453_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_453_inst_req_1;
      type_cast_453_inst_ack_1<= rack(0);
      type_cast_453_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_453_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call68_450,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_454,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_466_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_466_inst_req_0;
      type_cast_466_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_466_inst_req_1;
      type_cast_466_inst_ack_1<= rack(0);
      type_cast_466_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_466_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call73_463,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_467,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_478_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_478_inst_req_0;
      type_cast_478_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_478_inst_req_1;
      type_cast_478_inst_ack_1<= rack(0);
      type_cast_478_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_478_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call77_475,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv80_479,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_491_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_491_inst_req_0;
      type_cast_491_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_491_inst_req_1;
      type_cast_491_inst_ack_1<= rack(0);
      type_cast_491_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_491_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call82_488,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_492,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_503_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_503_inst_req_0;
      type_cast_503_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_503_inst_req_1;
      type_cast_503_inst_ack_1<= rack(0);
      type_cast_503_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_503_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call86_500,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv89_504,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_516_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_516_inst_req_0;
      type_cast_516_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_516_inst_req_1;
      type_cast_516_inst_ack_1<= rack(0);
      type_cast_516_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_516_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call91_513,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv92_517,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_528_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_528_inst_req_0;
      type_cast_528_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_528_inst_req_1;
      type_cast_528_inst_ack_1<= rack(0);
      type_cast_528_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_528_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call98_525,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv101_529,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_541_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_541_inst_req_0;
      type_cast_541_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_541_inst_req_1;
      type_cast_541_inst_ack_1<= rack(0);
      type_cast_541_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_541_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call103_538,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_542,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_553_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_553_inst_req_0;
      type_cast_553_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_553_inst_req_1;
      type_cast_553_inst_ack_1<= rack(0);
      type_cast_553_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_553_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call107_550,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv110_554,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_566_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_566_inst_req_0;
      type_cast_566_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_566_inst_req_1;
      type_cast_566_inst_ack_1<= rack(0);
      type_cast_566_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_566_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call112_563,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_567,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_578_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_578_inst_req_0;
      type_cast_578_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_578_inst_req_1;
      type_cast_578_inst_ack_1<= rack(0);
      type_cast_578_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_578_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call116_575,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv119_579,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_591_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_591_inst_req_0;
      type_cast_591_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_591_inst_req_1;
      type_cast_591_inst_ack_1<= rack(0);
      type_cast_591_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_591_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call121_588,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv122_592,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_601_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_601_inst_req_0;
      type_cast_601_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_601_inst_req_1;
      type_cast_601_inst_ack_1<= rack(0);
      type_cast_601_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_601_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_297,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv128_602,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_605_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_605_inst_req_0;
      type_cast_605_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_605_inst_req_1;
      type_cast_605_inst_ack_1<= rack(0);
      type_cast_605_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_605_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_347,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv130_606,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_609_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_609_inst_req_0;
      type_cast_609_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_609_inst_req_1;
      type_cast_609_inst_ack_1<= rack(0);
      type_cast_609_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_609_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add43_397,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv132_610,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_623_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_623_inst_req_0;
      type_cast_623_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_623_inst_req_1;
      type_cast_623_inst_ack_1<= rack(0);
      type_cast_623_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_623_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add33_372,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv138_624,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_627_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_627_inst_req_0;
      type_cast_627_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_627_inst_req_1;
      type_cast_627_inst_ack_1<= rack(0);
      type_cast_627_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_627_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_422,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv141_628,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_641_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_641_inst_req_0;
      type_cast_641_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_641_inst_req_1;
      type_cast_641_inst_ack_1<= rack(0);
      type_cast_641_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_641_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add75_472,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv147_642,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_645_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_645_inst_req_0;
      type_cast_645_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_645_inst_req_1;
      type_cast_645_inst_ack_1<= rack(0);
      type_cast_645_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_645_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add84_497,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv150_646,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_695_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_695_inst_req_0;
      type_cast_695_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_695_inst_req_1;
      type_cast_695_inst_ack_1<= rack(0);
      type_cast_695_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_695_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp409x_xop_692,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_27_696,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_718_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_718_inst_req_0;
      type_cast_718_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_718_inst_req_1;
      type_cast_718_inst_ack_1<= rack(0);
      type_cast_718_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_718_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext403_869,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_718_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_732_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_732_inst_req_0;
      type_cast_732_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_732_inst_req_1;
      type_cast_732_inst_ack_1<= rack(0);
      type_cast_732_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_732_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call160_729,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv161_733,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_745_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_745_inst_req_0;
      type_cast_745_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_745_inst_req_1;
      type_cast_745_inst_ack_1<= rack(0);
      type_cast_745_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_745_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call164_742,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv166_746,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_763_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_763_inst_req_0;
      type_cast_763_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_763_inst_req_1;
      type_cast_763_inst_ack_1<= rack(0);
      type_cast_763_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_763_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call170_760,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv172_764,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_781_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_781_inst_req_0;
      type_cast_781_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_781_inst_req_1;
      type_cast_781_inst_ack_1<= rack(0);
      type_cast_781_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_781_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call176_778,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv178_782,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_799_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_799_inst_req_0;
      type_cast_799_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_799_inst_req_1;
      type_cast_799_inst_ack_1<= rack(0);
      type_cast_799_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_799_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call182_796,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv184_800,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_817_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_817_inst_req_0;
      type_cast_817_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_817_inst_req_1;
      type_cast_817_inst_ack_1<= rack(0);
      type_cast_817_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_817_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call188_814,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv190_818,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_835_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_835_inst_req_0;
      type_cast_835_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_835_inst_req_1;
      type_cast_835_inst_ack_1<= rack(0);
      type_cast_835_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_835_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call194_832,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv196_836,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_853_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_853_inst_req_0;
      type_cast_853_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_853_inst_req_1;
      type_cast_853_inst_ack_1<= rack(0);
      type_cast_853_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_853_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call200_850,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv202_854,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_933_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_933_inst_req_0;
      type_cast_933_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_933_inst_req_1;
      type_cast_933_inst_ack_1<= rack(0);
      type_cast_933_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_933_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp395x_xop_930,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_40_934,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_956_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_956_inst_req_0;
      type_cast_956_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_956_inst_req_1;
      type_cast_956_inst_ack_1<= rack(0);
      type_cast_956_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_956_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext389_965,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_956_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1043_index_1_rename
    process(R_indvar_1042_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1042_resized;
      ov(13 downto 0) := iv;
      R_indvar_1042_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1043_index_1_resize
    process(indvar_1031) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1031;
      ov := iv(13 downto 0);
      R_indvar_1042_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1043_root_address_inst
    process(array_obj_ref_1043_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1043_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1043_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1194_index_1_rename
    process(R_shr307364_1193_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_shr307364_1193_resized;
      ov(13 downto 0) := iv;
      R_shr307364_1193_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1194_index_1_resize
    process(shr307364_1189) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shr307364_1189;
      ov := iv(13 downto 0);
      R_shr307364_1193_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1194_root_address_inst
    process(array_obj_ref_1194_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1194_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1194_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1215_index_1_rename
    process(R_shr313366_1214_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_shr313366_1214_resized;
      ov(13 downto 0) := iv;
      R_shr313366_1214_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1215_index_1_resize
    process(shr313366_1210) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shr313366_1210;
      ov := iv(13 downto 0);
      R_shr313366_1214_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1215_root_address_inst
    process(array_obj_ref_1215_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1215_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1215_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_724_index_1_rename
    process(R_indvar402_723_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar402_723_resized;
      ov(13 downto 0) := iv;
      R_indvar402_723_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_724_index_1_resize
    process(indvar402_712) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar402_712;
      ov := iv(13 downto 0);
      R_indvar402_723_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_724_root_address_inst
    process(array_obj_ref_724_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_724_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_724_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1047_addr_0
    process(ptr_deref_1047_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1047_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1047_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1047_base_resize
    process(arrayidx231_1045) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx231_1045;
      ov := iv(13 downto 0);
      ptr_deref_1047_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1047_gather_scatter
    process(type_cast_1049_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1049_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1047_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1047_root_address_inst
    process(ptr_deref_1047_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1047_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1047_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1199_addr_0
    process(ptr_deref_1199_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1199_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1199_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1199_base_resize
    process(arrayidx309_1196) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx309_1196;
      ov := iv(13 downto 0);
      ptr_deref_1199_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1199_gather_scatter
    process(ptr_deref_1199_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1199_data_0;
      ov(63 downto 0) := iv;
      tmp310_1200 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1199_root_address_inst
    process(ptr_deref_1199_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1199_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1199_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1219_addr_0
    process(ptr_deref_1219_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1219_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1219_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1219_base_resize
    process(arrayidx315_1217) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx315_1217;
      ov := iv(13 downto 0);
      ptr_deref_1219_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1219_gather_scatter
    process(tmp310_1200) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp310_1200;
      ov(63 downto 0) := iv;
      ptr_deref_1219_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1219_root_address_inst
    process(ptr_deref_1219_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1219_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1219_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_861_addr_0
    process(ptr_deref_861_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_861_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_861_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_861_base_resize
    process(arrayidx_726) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_726;
      ov := iv(13 downto 0);
      ptr_deref_861_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_861_gather_scatter
    process(add203_859) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add203_859;
      ov(63 downto 0) := iv;
      ptr_deref_861_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_861_root_address_inst
    process(ptr_deref_861_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_861_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_861_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1062_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1061;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1062_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1062_branch_req_0,
          ack0 => if_stmt_1062_branch_ack_0,
          ack1 => if_stmt_1062_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1275_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp342_1274;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1275_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1275_branch_req_0,
          ack0 => if_stmt_1275_branch_ack_0,
          ack1 => if_stmt_1275_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_668_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp376_667;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_668_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_668_branch_req_0,
          ack0 => if_stmt_668_branch_ack_0,
          ack1 => if_stmt_668_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_875_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_874;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_875_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_875_branch_req_0,
          ack0 => if_stmt_875_branch_ack_0,
          ack1 => if_stmt_875_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_891_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp212372_890;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_891_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_891_branch_req_0,
          ack0 => if_stmt_891_branch_ack_0,
          ack1 => if_stmt_891_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_971_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_970;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_971_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_971_branch_req_0,
          ack0 => if_stmt_971_branch_ack_0,
          ack1 => if_stmt_971_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_987_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp226369_986;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_987_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_987_branch_req_0,
          ack0 => if_stmt_987_branch_ack_0,
          ack1 => if_stmt_987_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1078_inst
    process(add75_472) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add75_472, type_cast_1077_wire_constant, tmp_var);
      add257_1079 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1089_inst
    process(add84_497) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add84_497, type_cast_1088_wire_constant, tmp_var);
      add269_1090 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1128_inst
    process(sub_1084, mul254_1124) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1084, mul254_1124, tmp_var);
      sub260_1129 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1143_inst
    process(input_dim1x_x1_1105, mul285_1139) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1105, mul285_1139, tmp_var);
      add286_1144 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1153_inst
    process(mul287_1149, input_dim2x_x0_1112) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul287_1149, input_dim2x_x0_1112, tmp_var);
      add288_1154 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1163_inst
    process(sub272_1095, mul266_1134) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub272_1095, mul266_1134, tmp_var);
      sub273_1164 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1168_inst
    process(sub273_1164, mul300_1159) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub273_1164, mul300_1159, tmp_var);
      add301_1169 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1178_inst
    process(mul302_1174, input_dim2x_x0_1112) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul302_1174, input_dim2x_x0_1112, tmp_var);
      add303_1179 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1226_inst
    process(input_dim2x_x0_1112) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x0_1112, type_cast_1225_wire_constant, tmp_var);
      add318_1227 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1240_inst
    process(inc327_1236, input_dim1x_x1_1105) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc327_1236, input_dim1x_x1_1105, tmp_var);
      inc327x_xinput_dim1x_x1_1241 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1261_inst
    process(inc336_1257, input_dim0x_x1_1098) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc336_1257, input_dim0x_x1_1098, tmp_var);
      inc336x_xinput_dim0x_x1_1262 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1010_inst
    process(tmp383_999) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp383_999, type_cast_1009_wire_constant, tmp_var);
      tmp383x_xop_1011 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_691_inst
    process(tmp409_680) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp409_680, type_cast_690_wire_constant, tmp_var);
      tmp409x_xop_692 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_929_inst
    process(tmp395_918) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp395_918, type_cast_928_wire_constant, tmp_var);
      tmp395x_xop_930 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1020_inst
    process(iNsTr_47_1015) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_47_1015, type_cast_1019_wire_constant, tmp_var);
      xx_xop_1021 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1055_inst
    process(indvar_1031) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1031, type_cast_1054_wire_constant, tmp_var);
      indvarx_xnext_1056 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_701_inst
    process(iNsTr_27_696) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_27_696, type_cast_700_wire_constant, tmp_var);
      xx_xop417_702 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_868_inst
    process(indvar402_712) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar402_712, type_cast_867_wire_constant, tmp_var);
      indvarx_xnext403_869 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_939_inst
    process(iNsTr_40_934) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_40_934, type_cast_938_wire_constant, tmp_var);
      xx_xop416_940 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_964_inst
    process(iNsTr_44_950) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_44_950, type_cast_963_wire_constant, tmp_var);
      indvarx_xnext389_965 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1231_inst
    process(add318_1227, add43_397) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(add318_1227, add43_397, tmp_var);
      cmp324_1232 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1252_inst
    process(inc327x_xinput_dim1x_x1_1241, add23_347) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc327x_xinput_dim1x_x1_1241, add23_347, tmp_var);
      cmp332_1253 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1273_inst
    process(inc336x_xinput_dim0x_x1_1262, add_297) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc336x_xinput_dim0x_x1_1262, add_297, tmp_var);
      cmp342_1274 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1060_inst
    process(indvarx_xnext_1056, tmp387_1028) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1056, tmp387_1028, tmp_var);
      exitcond1_1061 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_873_inst
    process(indvarx_xnext403_869, tmp414_709) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext403_869, tmp414_709, tmp_var);
      exitcond2_874 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_969_inst
    process(indvarx_xnext389_965, tmp400_947) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext389_965, tmp400_947, tmp_var);
      exitcond_970 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_679_inst
    process(mul133_620) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul133_620, type_cast_678_wire_constant, tmp_var);
      tmp409_680 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_917_inst
    process(tmp394_912) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp394_912, type_cast_916_wire_constant, tmp_var);
      tmp395_918 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_998_inst
    process(mul142_638) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul142_638, type_cast_997_wire_constant, tmp_var);
      tmp383_999 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1188_inst
    process(conv306_1183) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv306_1183, type_cast_1187_wire_constant, tmp_var);
      shr307364_1189 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1209_inst
    process(conv312_1204) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv312_1204, type_cast_1208_wire_constant, tmp_var);
      shr313366_1210 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1123_inst
    process(input_dim0x_x1_1098, add105_547) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x1_1098, add105_547, tmp_var);
      mul254_1124 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1133_inst
    process(input_dim1x_x1_1105, add114_572) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1105, add114_572, tmp_var);
      mul266_1134 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1138_inst
    process(input_dim0x_x1_1098, add23_347) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x1_1098, add23_347, tmp_var);
      mul285_1139 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1148_inst
    process(add286_1144, add43_397) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add286_1144, add43_397, tmp_var);
      mul287_1149 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1158_inst
    process(sub260_1129, add33_372) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub260_1129, add33_372, tmp_var);
      mul300_1159 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1173_inst
    process(add301_1169, add53_422) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add301_1169, add53_422, tmp_var);
      mul302_1174 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_614_inst
    process(conv130_606, conv128_602) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv130_606, conv128_602, tmp_var);
      mul_615 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_619_inst
    process(mul_615, conv132_610) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_615, conv132_610, tmp_var);
      mul133_620 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_632_inst
    process(conv138_624, add13_322) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv138_624, add13_322, tmp_var);
      mul139_633 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_637_inst
    process(mul139_633, conv141_628) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul139_633, conv141_628, tmp_var);
      mul142_638 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_650_inst
    process(conv147_642, add66_447) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv147_642, add66_447, tmp_var);
      mul148_651 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_655_inst
    process(mul148_651, conv150_646) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul148_651, conv150_646, tmp_var);
      mul151_656 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_660_inst
    process(mul151_656, add93_522) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul151_656, add93_522, tmp_var);
      mul154_661 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_901_inst
    process(add66_447, add93_522) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add66_447, add93_522, tmp_var);
      tmp390_902 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_906_inst
    process(tmp390_902, conv147_642) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp390_902, conv147_642, tmp_var);
      tmp392_907 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_911_inst
    process(tmp392_907, conv150_646) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp392_907, conv150_646, tmp_var);
      tmp394_912 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_296_inst
    process(shl_285, conv3_292) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_285, conv3_292, tmp_var);
      add_297 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_346_inst
    process(shl20_335, conv22_342) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl20_335, conv22_342, tmp_var);
      add23_347 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_371_inst
    process(shl30_360, conv32_367) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl30_360, conv32_367, tmp_var);
      add33_372 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_396_inst
    process(shl40_385, conv42_392) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl40_385, conv42_392, tmp_var);
      add43_397 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_421_inst
    process(shl50_410, conv52_417) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl50_410, conv52_417, tmp_var);
      add53_422 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_471_inst
    process(shl72_460, conv74_467) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl72_460, conv74_467, tmp_var);
      add75_472 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_496_inst
    process(shl81_485, conv83_492) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl81_485, conv83_492, tmp_var);
      add84_497 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_546_inst
    process(shl102_535, conv104_542) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl102_535, conv104_542, tmp_var);
      add105_547 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_571_inst
    process(shl111_560, conv113_567) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl111_560, conv113_567, tmp_var);
      add114_572 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_596_inst
    process(shl120_585, conv122_592) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl120_585, conv122_592, tmp_var);
      add123_597 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_321_inst
    process(shl10_310, conv12_317) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl10_310, conv12_317, tmp_var);
      add13_322 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_446_inst
    process(shl63_435, conv65_442) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl63_435, conv65_442, tmp_var);
      add66_447 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_521_inst
    process(shl90_510, conv92_517) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl90_510, conv92_517, tmp_var);
      add93_522 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_750_inst
    process(shl163_739, conv166_746) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl163_739, conv166_746, tmp_var);
      add167_751 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_768_inst
    process(shl169_757, conv172_764) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl169_757, conv172_764, tmp_var);
      add173_769 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_786_inst
    process(shl175_775, conv178_782) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl175_775, conv178_782, tmp_var);
      add179_787 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_804_inst
    process(shl181_793, conv184_800) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl181_793, conv184_800, tmp_var);
      add185_805 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_822_inst
    process(shl187_811, conv190_818) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl187_811, conv190_818, tmp_var);
      add191_823 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_840_inst
    process(shl193_829, conv196_836) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl193_829, conv196_836, tmp_var);
      add197_841 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_858_inst
    process(shl199_847, conv202_854) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl199_847, conv202_854, tmp_var);
      add203_859 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_284_inst
    process(conv1_279) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_279, type_cast_283_wire_constant, tmp_var);
      shl_285 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_334_inst
    process(conv19_329) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv19_329, type_cast_333_wire_constant, tmp_var);
      shl20_335 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_359_inst
    process(conv29_354) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv29_354, type_cast_358_wire_constant, tmp_var);
      shl30_360 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_384_inst
    process(conv39_379) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv39_379, type_cast_383_wire_constant, tmp_var);
      shl40_385 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_409_inst
    process(conv49_404) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv49_404, type_cast_408_wire_constant, tmp_var);
      shl50_410 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_459_inst
    process(conv71_454) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv71_454, type_cast_458_wire_constant, tmp_var);
      shl72_460 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_484_inst
    process(conv80_479) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv80_479, type_cast_483_wire_constant, tmp_var);
      shl81_485 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_534_inst
    process(conv101_529) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv101_529, type_cast_533_wire_constant, tmp_var);
      shl102_535 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_559_inst
    process(conv110_554) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv110_554, type_cast_558_wire_constant, tmp_var);
      shl111_560 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_584_inst
    process(conv119_579) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv119_579, type_cast_583_wire_constant, tmp_var);
      shl120_585 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_309_inst
    process(conv9_304) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv9_304, type_cast_308_wire_constant, tmp_var);
      shl10_310 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_434_inst
    process(conv62_429) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv62_429, type_cast_433_wire_constant, tmp_var);
      shl63_435 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_509_inst
    process(conv89_504) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv89_504, type_cast_508_wire_constant, tmp_var);
      shl90_510 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_738_inst
    process(conv161_733) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv161_733, type_cast_737_wire_constant, tmp_var);
      shl163_739 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_756_inst
    process(add167_751) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add167_751, type_cast_755_wire_constant, tmp_var);
      shl169_757 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_774_inst
    process(add173_769) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add173_769, type_cast_773_wire_constant, tmp_var);
      shl175_775 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_792_inst
    process(add179_787) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add179_787, type_cast_791_wire_constant, tmp_var);
      shl181_793 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_810_inst
    process(add185_805) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add185_805, type_cast_809_wire_constant, tmp_var);
      shl187_811 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_828_inst
    process(add191_823) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add191_823, type_cast_827_wire_constant, tmp_var);
      shl193_829 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_846_inst
    process(add197_841) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add197_841, type_cast_845_wire_constant, tmp_var);
      shl199_847 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1083_inst
    process(add257_1079, add123_597) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add257_1079, add123_597, tmp_var);
      sub_1084 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1094_inst
    process(add269_1090, add123_597) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add269_1090, add123_597, tmp_var);
      sub272_1095 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1299_inst
    process(conv349_1295, conv238_1287) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv349_1295, conv238_1287, tmp_var);
      sub353_1300 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1004_inst
    process(tmp383_999) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp383_999, type_cast_1003_wire_constant, tmp_var);
      tmp384_1005 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_666_inst
    process(mul133_620) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul133_620, type_cast_665_wire_constant, tmp_var);
      cmp376_667 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_685_inst
    process(tmp409_680) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp409_680, type_cast_684_wire_constant, tmp_var);
      tmp410_686 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_889_inst
    process(mul154_661) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul154_661, type_cast_888_wire_constant, tmp_var);
      cmp212372_890 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_923_inst
    process(tmp395_918) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp395_918, type_cast_922_wire_constant, tmp_var);
      tmp396_924 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_985_inst
    process(mul142_638) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul142_638, type_cast_984_wire_constant, tmp_var);
      cmp226369_986 <= tmp_var; --
    end process;
    -- shared split operator group (96) : array_obj_ref_1043_index_offset 
    ApIntAdd_group_96: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1042_scaled;
      array_obj_ref_1043_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1043_index_offset_req_0;
      array_obj_ref_1043_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1043_index_offset_req_1;
      array_obj_ref_1043_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_96_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_96_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_96",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 96
    -- shared split operator group (97) : array_obj_ref_1194_index_offset 
    ApIntAdd_group_97: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_shr307364_1193_scaled;
      array_obj_ref_1194_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1194_index_offset_req_0;
      array_obj_ref_1194_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1194_index_offset_req_1;
      array_obj_ref_1194_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_97_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_97_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_97",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 97
    -- shared split operator group (98) : array_obj_ref_1215_index_offset 
    ApIntAdd_group_98: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_shr313366_1214_scaled;
      array_obj_ref_1215_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1215_index_offset_req_0;
      array_obj_ref_1215_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1215_index_offset_req_1;
      array_obj_ref_1215_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_98_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_98_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_98",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 98
    -- shared split operator group (99) : array_obj_ref_724_index_offset 
    ApIntAdd_group_99: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar402_723_scaled;
      array_obj_ref_724_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_724_index_offset_req_0;
      array_obj_ref_724_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_724_index_offset_req_1;
      array_obj_ref_724_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_99_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_99_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_99",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 99
    -- unary operator type_cast_1285_inst
    process(call237_1072) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call237_1072, tmp_var);
      type_cast_1285_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1293_inst
    process(call348_1290) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call348_1290, tmp_var);
      type_cast_1293_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1199_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1199_load_0_req_0;
      ptr_deref_1199_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1199_load_0_req_1;
      ptr_deref_1199_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1199_word_address_0;
      ptr_deref_1199_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1047_store_0 ptr_deref_1219_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1047_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1219_store_0_req_0;
      ptr_deref_1047_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1219_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1047_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1219_store_0_req_1;
      ptr_deref_1047_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1219_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1047_word_address_0 & ptr_deref_1219_word_address_0;
      data_in <= ptr_deref_1047_data_0 & ptr_deref_1219_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_861_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_861_store_0_req_0;
      ptr_deref_861_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_861_store_0_req_1;
      ptr_deref_861_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_861_word_address_0;
      data_in <= ptr_deref_861_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared inport operator group (0) : RPIPE_ConvTranspose_input_pipe_273_inst RPIPE_ConvTranspose_input_pipe_287_inst RPIPE_ConvTranspose_input_pipe_299_inst RPIPE_ConvTranspose_input_pipe_312_inst RPIPE_ConvTranspose_input_pipe_324_inst RPIPE_ConvTranspose_input_pipe_337_inst RPIPE_ConvTranspose_input_pipe_349_inst RPIPE_ConvTranspose_input_pipe_362_inst RPIPE_ConvTranspose_input_pipe_374_inst RPIPE_ConvTranspose_input_pipe_387_inst RPIPE_ConvTranspose_input_pipe_399_inst RPIPE_ConvTranspose_input_pipe_412_inst RPIPE_ConvTranspose_input_pipe_424_inst RPIPE_ConvTranspose_input_pipe_437_inst RPIPE_ConvTranspose_input_pipe_449_inst RPIPE_ConvTranspose_input_pipe_462_inst RPIPE_ConvTranspose_input_pipe_474_inst RPIPE_ConvTranspose_input_pipe_487_inst RPIPE_ConvTranspose_input_pipe_499_inst RPIPE_ConvTranspose_input_pipe_512_inst RPIPE_ConvTranspose_input_pipe_524_inst RPIPE_ConvTranspose_input_pipe_537_inst RPIPE_ConvTranspose_input_pipe_549_inst RPIPE_ConvTranspose_input_pipe_562_inst RPIPE_ConvTranspose_input_pipe_574_inst RPIPE_ConvTranspose_input_pipe_587_inst RPIPE_ConvTranspose_input_pipe_728_inst RPIPE_ConvTranspose_input_pipe_741_inst RPIPE_ConvTranspose_input_pipe_759_inst RPIPE_ConvTranspose_input_pipe_777_inst RPIPE_ConvTranspose_input_pipe_795_inst RPIPE_ConvTranspose_input_pipe_813_inst RPIPE_ConvTranspose_input_pipe_831_inst RPIPE_ConvTranspose_input_pipe_849_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(271 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 33 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 33 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 33 downto 0);
      signal guard_vector : std_logic_vector( 33 downto 0);
      constant outBUFs : IntegerArray(33 downto 0) := (33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(33 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false);
      constant guardBuffering: IntegerArray(33 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2);
      -- 
    begin -- 
      reqL_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_273_inst_req_0;
      reqL_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_287_inst_req_0;
      reqL_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_299_inst_req_0;
      reqL_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_312_inst_req_0;
      reqL_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_324_inst_req_0;
      reqL_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_337_inst_req_0;
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_349_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_362_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_374_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_387_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_399_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_412_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_424_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_437_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_449_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_462_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_474_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_487_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_499_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_512_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_524_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_537_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_549_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_562_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_574_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_587_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_728_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_741_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_759_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_777_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_795_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_813_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_831_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_849_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_273_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_287_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_299_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_312_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_324_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_337_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_349_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_362_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_374_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_387_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_399_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_412_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_424_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_437_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_449_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_462_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_474_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_487_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_499_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_512_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_524_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_537_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_549_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_562_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_574_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_587_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_728_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_741_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_759_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_777_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_795_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_813_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_831_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_849_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_273_inst_req_1;
      reqR_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_287_inst_req_1;
      reqR_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_299_inst_req_1;
      reqR_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_312_inst_req_1;
      reqR_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_324_inst_req_1;
      reqR_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_337_inst_req_1;
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_349_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_362_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_374_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_387_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_399_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_412_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_424_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_437_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_449_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_462_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_474_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_487_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_499_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_512_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_524_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_537_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_549_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_562_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_574_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_587_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_728_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_741_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_759_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_777_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_795_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_813_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_831_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_849_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_273_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_287_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_299_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_312_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_324_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_337_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_349_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_362_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_374_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_387_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_399_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_412_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_424_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_437_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_449_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_462_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_474_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_487_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_499_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_512_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_524_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_537_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_549_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_562_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_574_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_587_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_728_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_741_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_759_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_777_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_795_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_813_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_831_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_849_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      call_274 <= data_out(271 downto 264);
      call2_288 <= data_out(263 downto 256);
      call6_300 <= data_out(255 downto 248);
      call11_313 <= data_out(247 downto 240);
      call16_325 <= data_out(239 downto 232);
      call21_338 <= data_out(231 downto 224);
      call26_350 <= data_out(223 downto 216);
      call31_363 <= data_out(215 downto 208);
      call36_375 <= data_out(207 downto 200);
      call41_388 <= data_out(199 downto 192);
      call46_400 <= data_out(191 downto 184);
      call51_413 <= data_out(183 downto 176);
      call59_425 <= data_out(175 downto 168);
      call64_438 <= data_out(167 downto 160);
      call68_450 <= data_out(159 downto 152);
      call73_463 <= data_out(151 downto 144);
      call77_475 <= data_out(143 downto 136);
      call82_488 <= data_out(135 downto 128);
      call86_500 <= data_out(127 downto 120);
      call91_513 <= data_out(119 downto 112);
      call98_525 <= data_out(111 downto 104);
      call103_538 <= data_out(103 downto 96);
      call107_550 <= data_out(95 downto 88);
      call112_563 <= data_out(87 downto 80);
      call116_575 <= data_out(79 downto 72);
      call121_588 <= data_out(71 downto 64);
      call160_729 <= data_out(63 downto 56);
      call164_742 <= data_out(55 downto 48);
      call170_760 <= data_out(47 downto 40);
      call176_778 <= data_out(39 downto 32);
      call182_796 <= data_out(31 downto 24);
      call188_814 <= data_out(23 downto 16);
      call194_832 <= data_out(15 downto 8);
      call200_850 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_0_gI", nreqs => 34, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_0", data_width => 8,  num_reqs => 34,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_elapsed_time_pipe_1301_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1301_inst_req_0;
      WPIPE_elapsed_time_pipe_1301_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1301_inst_req_1;
      WPIPE_elapsed_time_pipe_1301_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub353_1300;
      elapsed_time_pipe_write_0_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1072_call call_stmt_1290_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1072_call_req_0;
      reqL_unguarded(0) <= call_stmt_1290_call_req_0;
      call_stmt_1072_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1290_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1072_call_req_1;
      reqR_unguarded(0) <= call_stmt_1290_call_req_1;
      call_stmt_1072_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1290_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call237_1072 <= data_out(127 downto 64);
      call348_1290 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1306_call 
    sendOutput_call_group_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1306_call_req_0;
      call_stmt_1306_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1306_call_req_1;
      call_stmt_1306_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendOutput_call_group_1_gI: SplitGuardInterface generic map(name => "sendOutput_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= mul142_638;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 32,
        owidth => 32,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => sendOutput_call_reqs(0),
          ackR => sendOutput_call_acks(0),
          dataR => sendOutput_call_data(31 downto 0),
          tagR => sendOutput_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendOutput_return_acks(0), -- cross-over
          ackL => sendOutput_return_reqs(0), -- cross-over
          tagL => sendOutput_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_959_call 
    fill_kernel_call_group_2: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_959_call_req_0;
      call_stmt_959_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_959_call_req_1;
      call_stmt_959_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      fill_kernel_call_group_2_gI: SplitGuardInterface generic map(name => "fill_kernel_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= iNsTr_44_950;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 64,
        owidth => 64,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => fill_kernel_call_reqs(0),
          ackR => fill_kernel_call_acks(0),
          dataR => fill_kernel_call_data(63 downto 0),
          tagR => fill_kernel_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => fill_kernel_return_acks(0), -- cross-over
          ackL => fill_kernel_return_reqs(0), -- cross-over
          tagL => fill_kernel_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity fill_kernel is -- 
  generic (tag_length : integer); 
  port ( -- 
    addr : in  std_logic_vector(63 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(11 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity fill_kernel;
architecture fill_kernel_arch of fill_kernel is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal addr_buffer :  std_logic_vector(63 downto 0);
  signal addr_update_enable: Boolean;
  -- output port buffer signals
  signal fill_kernel_CP_0_start: Boolean;
  signal fill_kernel_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal CONCAT_u48_u64_47_inst_req_1 : boolean;
  signal CONCAT_u48_u64_47_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_39_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_39_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_39_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_39_inst_ack_1 : boolean;
  signal CONCAT_u8_u16_40_inst_req_0 : boolean;
  signal CONCAT_u8_u16_40_inst_ack_0 : boolean;
  signal CONCAT_u8_u16_40_inst_req_1 : boolean;
  signal CONCAT_u8_u16_40_inst_ack_1 : boolean;
  signal CONCAT_u48_u64_47_inst_req_0 : boolean;
  signal CONCAT_u48_u64_47_inst_ack_0 : boolean;
  signal array_obj_ref_62_index_offset_req_0 : boolean;
  signal array_obj_ref_62_index_offset_ack_0 : boolean;
  signal array_obj_ref_62_index_offset_req_1 : boolean;
  signal if_stmt_49_branch_req_0 : boolean;
  signal if_stmt_49_branch_ack_1 : boolean;
  signal if_stmt_49_branch_ack_0 : boolean;
  signal phi_stmt_23_req_0 : boolean;
  signal phi_stmt_17_req_0 : boolean;
  signal ninput_word_48_27_buf_req_0 : boolean;
  signal ninput_word_48_27_buf_ack_0 : boolean;
  signal ninput_word_48_27_buf_req_1 : boolean;
  signal ninput_word_48_27_buf_ack_1 : boolean;
  signal phi_stmt_23_req_1 : boolean;
  signal nmycount_33_22_buf_req_0 : boolean;
  signal nmycount_33_22_buf_ack_0 : boolean;
  signal nmycount_33_22_buf_req_1 : boolean;
  signal nmycount_33_22_buf_ack_1 : boolean;
  signal phi_stmt_17_req_1 : boolean;
  signal phi_stmt_17_ack_0 : boolean;
  signal phi_stmt_23_ack_0 : boolean;
  signal array_obj_ref_62_index_offset_ack_1 : boolean;
  signal addr_of_63_final_reg_req_0 : boolean;
  signal addr_of_63_final_reg_ack_0 : boolean;
  signal addr_of_63_final_reg_req_1 : boolean;
  signal addr_of_63_final_reg_ack_1 : boolean;
  signal ptr_deref_66_store_0_req_0 : boolean;
  signal ptr_deref_66_store_0_ack_0 : boolean;
  signal ptr_deref_66_store_0_req_1 : boolean;
  signal ptr_deref_66_store_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "fill_kernel_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 64) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= addr;
  addr_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(tag_length + 63 downto 64) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 63 downto 64);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  fill_kernel_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "fill_kernel_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= fill_kernel_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= fill_kernel_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= fill_kernel_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  fill_kernel_CP_0: Block -- control-path 
    signal fill_kernel_CP_0_elements: BooleanArray(33 downto 0);
    -- 
  begin -- 
    fill_kernel_CP_0_elements(0) <= fill_kernel_CP_0_start;
    fill_kernel_CP_0_symbol <= fill_kernel_CP_0_elements(33);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	12 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_15/$entry
      -- CP-element group 0: 	 branch_block_stmt_15/branch_block_stmt_15__entry__
      -- CP-element group 0: 	 branch_block_stmt_15/merge_stmt_16__entry__
      -- CP-element group 0: 	 branch_block_stmt_15/merge_stmt_16_dead_link/$entry
      -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	26 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	7 
    -- CP-element group 1: 	9 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (12) 
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_35_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u48_u64_47_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_35_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_35_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_15/merge_stmt_16__exit__
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48__entry__
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/$entry
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_update_start_
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u48_u64_47_update_start_
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u48_u64_47_Update/$entry
      -- 
    cr_71_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_71_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(1), ack => CONCAT_u48_u64_47_inst_req_1); -- 
    rr_24_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_24_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(1), ack => RPIPE_ConvTranspose_input_pipe_35_inst_req_0); -- 
    cr_57_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_57_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(1), ack => CONCAT_u8_u16_40_inst_req_1); -- 
    fill_kernel_CP_0_elements(1) <= fill_kernel_CP_0_elements(26);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_35_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_35_update_start_
      -- CP-element group 2: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_35_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_35_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_35_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_35_Update/cr
      -- 
    ra_25_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_35_inst_ack_0, ack => fill_kernel_CP_0_elements(2)); -- 
    cr_29_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_29_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(2), ack => RPIPE_ConvTranspose_input_pipe_35_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_35_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_35_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_35_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_39_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_39_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_39_Sample/rr
      -- 
    ca_30_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_35_inst_ack_1, ack => fill_kernel_CP_0_elements(3)); -- 
    rr_42_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_42_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(3), ack => RPIPE_ConvTranspose_input_pipe_39_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_39_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_39_update_start_
      -- CP-element group 4: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_39_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_39_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_39_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_39_Update/cr
      -- 
    ra_43_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_39_inst_ack_0, ack => fill_kernel_CP_0_elements(4)); -- 
    cr_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(4), ack => RPIPE_ConvTranspose_input_pipe_39_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_39_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_39_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_ConvTranspose_input_pipe_39_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_Sample/rr
      -- 
    ca_48_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_39_inst_ack_1, ack => fill_kernel_CP_0_elements(5)); -- 
    rr_52_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_52_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(5), ack => CONCAT_u8_u16_40_inst_req_0); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_Sample/ra
      -- 
    ra_53_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u8_u16_40_inst_ack_0, ack => fill_kernel_CP_0_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	1 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u48_u64_47_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u48_u64_47_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u48_u64_47_Sample/rr
      -- 
    ca_58_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u8_u16_40_inst_ack_1, ack => fill_kernel_CP_0_elements(7)); -- 
    rr_66_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_66_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(7), ack => CONCAT_u48_u64_47_inst_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u48_u64_47_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u48_u64_47_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u48_u64_47_Sample/ra
      -- 
    ra_67_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u48_u64_47_inst_ack_0, ack => fill_kernel_CP_0_elements(8)); -- 
    -- CP-element group 9:  branch  transition  place  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (27) 
      -- CP-element group 9: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u48_u64_47_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48__exit__
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49__entry__
      -- CP-element group 9: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/$exit
      -- CP-element group 9: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u48_u64_47_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u48_u64_47_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_dead_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/$entry
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/$exit
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/$entry
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/$exit
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/ULT_u4_u1_52_inputs/$entry
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/ULT_u4_u1_52_inputs/$exit
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/SplitProtocol/$entry
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/SplitProtocol/$exit
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/SplitProtocol/Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/SplitProtocol/Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/SplitProtocol/Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/SplitProtocol/Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/SplitProtocol/Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/SplitProtocol/Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/SplitProtocol/Update/cr
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/SplitProtocol/Update/ca
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/branch_req
      -- CP-element group 9: 	 branch_block_stmt_15/ULT_u4_u1_52_place
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_if_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_else_link/$entry
      -- 
    ca_72_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u48_u64_47_inst_ack_1, ack => fill_kernel_CP_0_elements(9)); -- 
    branch_req_99_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_99_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(9), ack => if_stmt_49_branch_req_0); -- 
    -- CP-element group 10:  fork  transition  place  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	16 
    -- CP-element group 10: 	17 
    -- CP-element group 10: 	19 
    -- CP-element group 10: 	20 
    -- CP-element group 10:  members (18) 
      -- CP-element group 10: 	 branch_block_stmt_15/if_stmt_49_if_link/$exit
      -- CP-element group 10: 	 branch_block_stmt_15/if_stmt_49_if_link/if_choice_transition
      -- CP-element group 10: 	 branch_block_stmt_15/loopback
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Sample/req
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Update/req
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Sample/req
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Update/req
      -- 
    if_choice_transition_104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_49_branch_ack_1, ack => fill_kernel_CP_0_elements(10)); -- 
    req_148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(10), ack => ninput_word_48_27_buf_req_0); -- 
    req_153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(10), ack => ninput_word_48_27_buf_req_1); -- 
    req_168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(10), ack => nmycount_33_22_buf_req_0); -- 
    req_173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(10), ack => nmycount_33_22_buf_req_1); -- 
    -- CP-element group 11:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	27 
    -- CP-element group 11: 	28 
    -- CP-element group 11: 	30 
    -- CP-element group 11: 	32 
    -- CP-element group 11:  members (30) 
      -- CP-element group 11: 	 branch_block_stmt_15/$exit
      -- CP-element group 11: 	 branch_block_stmt_15/branch_block_stmt_15__exit__
      -- CP-element group 11: 	 branch_block_stmt_15/if_stmt_49__exit__
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_update_start
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Sample/$entry
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Sample/req
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Update/$entry
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Update/req
      -- CP-element group 11: 	 branch_block_stmt_15/if_stmt_49_else_link/$exit
      -- CP-element group 11: 	 branch_block_stmt_15/if_stmt_49_else_link/else_choice_transition
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/$entry
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_update_start_
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_resized_1
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_scaled_1
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_computed_1
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_resize_1/$entry
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_resize_1/$exit
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_resize_1/index_resize_req
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_resize_1/index_resize_ack
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_scale_1/$entry
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_scale_1/$exit
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_scale_1/scale_rename_req
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_scale_1/scale_rename_ack
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_complete/$entry
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_complete/req
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_update_start_
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/$entry
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/word_access_complete/$entry
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/word_access_complete/word_0/$entry
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/word_access_complete/word_0/cr
      -- 
    else_choice_transition_108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_49_branch_ack_0, ack => fill_kernel_CP_0_elements(11)); -- 
    req_209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(11), ack => array_obj_ref_62_index_offset_req_0); -- 
    req_214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(11), ack => array_obj_ref_62_index_offset_req_1); -- 
    req_229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(11), ack => addr_of_63_final_reg_req_1); -- 
    cr_279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(11), ack => ptr_deref_66_store_0_req_1); -- 
    -- CP-element group 12:  fork  transition  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/$entry
      -- CP-element group 12: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_23/$entry
      -- CP-element group 12: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_23/phi_stmt_23_sources/$entry
      -- CP-element group 12: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_17/$entry
      -- CP-element group 12: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_17/phi_stmt_17_sources/$entry
      -- 
    fill_kernel_CP_0_elements(12) <= fill_kernel_CP_0_elements(0);
    -- CP-element group 13:  transition  output  delay-element  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (4) 
      -- CP-element group 13: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_23/$exit
      -- CP-element group 13: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_23/phi_stmt_23_sources/$exit
      -- CP-element group 13: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_23/phi_stmt_23_sources/type_cast_26_konst_delay_trans
      -- CP-element group 13: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_23/phi_stmt_23_req
      -- 
    phi_stmt_23_req_124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_23_req_124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(13), ack => phi_stmt_23_req_0); -- 
    -- Element group fill_kernel_CP_0_elements(13) is a control-delay.
    cp_element_13_delay: control_delay_element  generic map(name => " 13_delay", delay_value => 1)  port map(req => fill_kernel_CP_0_elements(12), ack => fill_kernel_CP_0_elements(13), clk => clk, reset =>reset);
    -- CP-element group 14:  transition  output  delay-element  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (4) 
      -- CP-element group 14: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_17/$exit
      -- CP-element group 14: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_17/phi_stmt_17_sources/$exit
      -- CP-element group 14: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_17/phi_stmt_17_sources/type_cast_21_konst_delay_trans
      -- CP-element group 14: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_17/phi_stmt_17_req
      -- 
    phi_stmt_17_req_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_17_req_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(14), ack => phi_stmt_17_req_0); -- 
    -- Element group fill_kernel_CP_0_elements(14) is a control-delay.
    cp_element_14_delay: control_delay_element  generic map(name => " 14_delay", delay_value => 1)  port map(req => fill_kernel_CP_0_elements(12), ack => fill_kernel_CP_0_elements(14), clk => clk, reset =>reset);
    -- CP-element group 15:  join  transition  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	23 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/$exit
      -- 
    fill_kernel_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "fill_kernel_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_kernel_CP_0_elements(13) & fill_kernel_CP_0_elements(14);
      gj_fill_kernel_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_kernel_CP_0_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	10 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Sample/ack
      -- 
    ack_149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ninput_word_48_27_buf_ack_0, ack => fill_kernel_CP_0_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	10 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Update/ack
      -- 
    ack_154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ninput_word_48_27_buf_ack_1, ack => fill_kernel_CP_0_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	22 
    -- CP-element group 18:  members (4) 
      -- CP-element group 18: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/$exit
      -- CP-element group 18: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/$exit
      -- CP-element group 18: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/$exit
      -- CP-element group 18: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_req
      -- 
    phi_stmt_23_req_155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_23_req_155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(18), ack => phi_stmt_23_req_1); -- 
    fill_kernel_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "fill_kernel_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_kernel_CP_0_elements(16) & fill_kernel_CP_0_elements(17);
      gj_fill_kernel_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_kernel_CP_0_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	10 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Sample/ack
      -- 
    ack_169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_33_22_buf_ack_0, ack => fill_kernel_CP_0_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	10 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Update/ack
      -- 
    ack_174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_33_22_buf_ack_1, ack => fill_kernel_CP_0_elements(20)); -- 
    -- CP-element group 21:  join  transition  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/$exit
      -- CP-element group 21: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/$exit
      -- CP-element group 21: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/$exit
      -- CP-element group 21: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_req
      -- 
    phi_stmt_17_req_175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_17_req_175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(21), ack => phi_stmt_17_req_1); -- 
    fill_kernel_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "fill_kernel_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_kernel_CP_0_elements(19) & fill_kernel_CP_0_elements(20);
      gj_fill_kernel_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_kernel_CP_0_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	18 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_15/loopback_PhiReq/$exit
      -- 
    fill_kernel_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "fill_kernel_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_kernel_CP_0_elements(18) & fill_kernel_CP_0_elements(21);
      gj_fill_kernel_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_kernel_CP_0_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  merge  fork  transition  place  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	15 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_15/merge_stmt_16_PhiReqMerge
      -- CP-element group 23: 	 branch_block_stmt_15/merge_stmt_16_PhiAck/$entry
      -- 
    fill_kernel_CP_0_elements(23) <= OrReduce(fill_kernel_CP_0_elements(15) & fill_kernel_CP_0_elements(22));
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_15/merge_stmt_16_PhiAck/phi_stmt_17_ack
      -- 
    phi_stmt_17_ack_180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_17_ack_0, ack => fill_kernel_CP_0_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_15/merge_stmt_16_PhiAck/phi_stmt_23_ack
      -- 
    phi_stmt_23_ack_181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_23_ack_0, ack => fill_kernel_CP_0_elements(25)); -- 
    -- CP-element group 26:  join  transition  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	1 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_15/merge_stmt_16_PhiAck/$exit
      -- 
    fill_kernel_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "fill_kernel_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_kernel_CP_0_elements(24) & fill_kernel_CP_0_elements(25);
      gj_fill_kernel_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_kernel_CP_0_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	11 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	33 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Sample/$exit
      -- CP-element group 27: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Sample/ack
      -- CP-element group 27: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_sample_complete
      -- 
    ack_210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_62_index_offset_ack_0, ack => fill_kernel_CP_0_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	11 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (11) 
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Update/$exit
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_sample_start_
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_root_address_calculated
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_offset_calculated
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Update/ack
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_base_plus_offset/$entry
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_base_plus_offset/$exit
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_base_plus_offset/sum_rename_req
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_base_plus_offset/sum_rename_ack
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_request/$entry
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_request/req
      -- 
    ack_215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_62_index_offset_ack_1, ack => fill_kernel_CP_0_elements(28)); -- 
    req_224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(28), ack => addr_of_63_final_reg_req_0); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_sample_completed_
      -- CP-element group 29: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_request/$exit
      -- CP-element group 29: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_request/ack
      -- 
    ack_225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_63_final_reg_ack_0, ack => fill_kernel_CP_0_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	11 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (28) 
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_update_completed_
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_complete/$exit
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_complete/ack
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_sample_start_
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_address_calculated
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_word_address_calculated
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_root_address_calculated
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_address_resized
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_addr_resize/$entry
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_addr_resize/$exit
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_addr_resize/base_resize_req
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_addr_resize/base_resize_ack
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_plus_offset/$entry
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_plus_offset/$exit
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_plus_offset/sum_rename_req
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_plus_offset/sum_rename_ack
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_word_addrgen/$entry
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_word_addrgen/$exit
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_word_addrgen/root_register_req
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_word_addrgen/root_register_ack
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/$entry
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/ptr_deref_66_Split/$entry
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/ptr_deref_66_Split/$exit
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/ptr_deref_66_Split/split_req
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/ptr_deref_66_Split/split_ack
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/word_access_start/$entry
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/word_access_start/word_0/$entry
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/word_access_start/word_0/rr
      -- 
    ack_230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_63_final_reg_ack_1, ack => fill_kernel_CP_0_elements(30)); -- 
    rr_268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_kernel_CP_0_elements(30), ack => ptr_deref_66_store_0_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_sample_completed_
      -- CP-element group 31: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/$exit
      -- CP-element group 31: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/word_access_start/$exit
      -- CP-element group 31: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/word_access_start/word_0/$exit
      -- CP-element group 31: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/word_access_start/word_0/ra
      -- 
    ra_269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_66_store_0_ack_0, ack => fill_kernel_CP_0_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	11 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_update_completed_
      -- CP-element group 32: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/$exit
      -- CP-element group 32: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/word_access_complete/$exit
      -- CP-element group 32: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/word_access_complete/word_0/$exit
      -- CP-element group 32: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/word_access_complete/word_0/ca
      -- 
    ca_280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_66_store_0_ack_1, ack => fill_kernel_CP_0_elements(32)); -- 
    -- CP-element group 33:  join  transition  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	27 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 $exit
      -- CP-element group 33: 	 assign_stmt_64_to_assign_stmt_68/$exit
      -- 
    fill_kernel_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "fill_kernel_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_kernel_CP_0_elements(27) & fill_kernel_CP_0_elements(32);
      gj_fill_kernel_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_kernel_CP_0_elements(33), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal RPIPE_ConvTranspose_input_pipe_39_wire : std_logic_vector(7 downto 0);
    signal R_addr_61_resized : std_logic_vector(11 downto 0);
    signal R_addr_61_scaled : std_logic_vector(11 downto 0);
    signal ULT_u4_u1_52_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_62_constant_part_of_offset : std_logic_vector(11 downto 0);
    signal array_obj_ref_62_final_offset : std_logic_vector(11 downto 0);
    signal array_obj_ref_62_offset_scale_factor_0 : std_logic_vector(11 downto 0);
    signal array_obj_ref_62_offset_scale_factor_1 : std_logic_vector(11 downto 0);
    signal array_obj_ref_62_resized_base_address : std_logic_vector(11 downto 0);
    signal array_obj_ref_62_root_address : std_logic_vector(11 downto 0);
    signal input_word_23 : std_logic_vector(63 downto 0);
    signal konst_31_wire_constant : std_logic_vector(3 downto 0);
    signal konst_51_wire_constant : std_logic_vector(3 downto 0);
    signal mycount_17 : std_logic_vector(3 downto 0);
    signal ninput_word_48 : std_logic_vector(63 downto 0);
    signal ninput_word_48_27_buffered : std_logic_vector(63 downto 0);
    signal nmycount_33 : std_logic_vector(3 downto 0);
    signal nmycount_33_22_buffered : std_logic_vector(3 downto 0);
    signal ptr_64 : std_logic_vector(31 downto 0);
    signal ptr_deref_66_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_66_resized_base_address : std_logic_vector(11 downto 0);
    signal ptr_deref_66_root_address : std_logic_vector(11 downto 0);
    signal ptr_deref_66_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_66_word_address_0 : std_logic_vector(11 downto 0);
    signal ptr_deref_66_word_offset_0 : std_logic_vector(11 downto 0);
    signal slice_45_wire : std_logic_vector(47 downto 0);
    signal type_cast_21_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_26_wire_constant : std_logic_vector(63 downto 0);
    signal val1_36 : std_logic_vector(7 downto 0);
    signal val_41 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_62_constant_part_of_offset <= "000000000000";
    array_obj_ref_62_offset_scale_factor_0 <= "000000000000";
    array_obj_ref_62_offset_scale_factor_1 <= "000000000001";
    array_obj_ref_62_resized_base_address <= "000000000000";
    konst_31_wire_constant <= "0001";
    konst_51_wire_constant <= "0011";
    ptr_deref_66_word_offset_0 <= "000000000000";
    type_cast_21_wire_constant <= "0000";
    type_cast_26_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_17: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_21_wire_constant & nmycount_33_22_buffered;
      req <= phi_stmt_17_req_0 & phi_stmt_17_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_17",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 4) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_17_ack_0,
          idata => idata,
          odata => mycount_17,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_17
    phi_stmt_23: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_26_wire_constant & ninput_word_48_27_buffered;
      req <= phi_stmt_23_req_0 & phi_stmt_23_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_23",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_23_ack_0,
          idata => idata,
          odata => input_word_23,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_23
    -- flow-through slice operator slice_45_inst
    slice_45_wire <= input_word_23(47 downto 0);
    addr_of_63_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_63_final_reg_req_0;
      addr_of_63_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_63_final_reg_req_1;
      addr_of_63_final_reg_ack_1<= rack(0);
      addr_of_63_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_63_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 12,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_62_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ptr_64,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    ninput_word_48_27_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= ninput_word_48_27_buf_req_0;
      ninput_word_48_27_buf_ack_0<= wack(0);
      rreq(0) <= ninput_word_48_27_buf_req_1;
      ninput_word_48_27_buf_ack_1<= rack(0);
      ninput_word_48_27_buf : InterlockBuffer generic map ( -- 
        name => "ninput_word_48_27_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ninput_word_48,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ninput_word_48_27_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_33_22_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_33_22_buf_req_0;
      nmycount_33_22_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_33_22_buf_req_1;
      nmycount_33_22_buf_ack_1<= rack(0);
      nmycount_33_22_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_33_22_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_33,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_33_22_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_62_index_1_rename
    process(R_addr_61_resized) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(11 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_61_resized;
      ov(11 downto 0) := iv;
      R_addr_61_scaled <= ov(11 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_62_index_1_resize
    process(addr_buffer) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(11 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_buffer;
      ov := iv(11 downto 0);
      R_addr_61_resized <= ov(11 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_62_root_address_inst
    process(array_obj_ref_62_final_offset) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(11 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_62_final_offset;
      ov(11 downto 0) := iv;
      array_obj_ref_62_root_address <= ov(11 downto 0);
      --
    end process;
    -- equivalence ptr_deref_66_addr_0
    process(ptr_deref_66_root_address) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(11 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_66_root_address;
      ov(11 downto 0) := iv;
      ptr_deref_66_word_address_0 <= ov(11 downto 0);
      --
    end process;
    -- equivalence ptr_deref_66_base_resize
    process(ptr_64) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(11 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_64;
      ov := iv(11 downto 0);
      ptr_deref_66_resized_base_address <= ov(11 downto 0);
      --
    end process;
    -- equivalence ptr_deref_66_gather_scatter
    process(ninput_word_48) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ninput_word_48;
      ov(63 downto 0) := iv;
      ptr_deref_66_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_66_root_address_inst
    process(ptr_deref_66_resized_base_address) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(11 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_66_resized_base_address;
      ov(11 downto 0) := iv;
      ptr_deref_66_root_address <= ov(11 downto 0);
      --
    end process;
    if_stmt_49_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u4_u1_52_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_49_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_49_branch_req_0,
          ack0 => if_stmt_49_branch_ack_0,
          ack1 => if_stmt_49_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u4_u4_32_inst
    process(mycount_17) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_17, konst_31_wire_constant, tmp_var);
      nmycount_33 <= tmp_var; --
    end process;
    -- shared split operator group (1) : CONCAT_u48_u64_47_inst 
    ApConcat_group_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= slice_45_wire & val_41;
      ninput_word_48 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u48_u64_47_inst_req_0;
      CONCAT_u48_u64_47_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u48_u64_47_inst_req_1;
      CONCAT_u48_u64_47_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_1_gI: SplitGuardInterface generic map(name => "ApConcat_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 48,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : CONCAT_u8_u16_40_inst 
    ApConcat_group_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= val1_36 & RPIPE_ConvTranspose_input_pipe_39_wire;
      val_41 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u8_u16_40_inst_req_0;
      CONCAT_u8_u16_40_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u8_u16_40_inst_req_1;
      CONCAT_u8_u16_40_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_2_gI: SplitGuardInterface generic map(name => "ApConcat_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- binary operator ULT_u4_u1_52_inst
    process(mycount_17) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_17, konst_51_wire_constant, tmp_var);
      ULT_u4_u1_52_wire <= tmp_var; --
    end process;
    -- shared split operator group (4) : array_obj_ref_62_index_offset 
    ApIntAdd_group_4: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr_61_scaled;
      array_obj_ref_62_final_offset <= data_out(11 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_62_index_offset_req_0;
      array_obj_ref_62_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_62_index_offset_req_1;
      array_obj_ref_62_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_4_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000000000000",
          constant_width => 12,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared store operator group (0) : ptr_deref_66_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(11 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_66_store_0_req_0;
      ptr_deref_66_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_66_store_0_req_1;
      ptr_deref_66_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_66_word_address_0;
      data_in <= ptr_deref_66_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 12,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(11 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_ConvTranspose_input_pipe_35_inst RPIPE_ConvTranspose_input_pipe_39_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_35_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_39_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_35_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_39_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_35_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_39_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_35_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_39_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      val1_36 <= data_out(15 downto 8);
      RPIPE_ConvTranspose_input_pipe_39_wire <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_0", data_width => 8,  num_reqs => 2,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end fill_kernel_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendOutput is -- 
  generic (tag_length : integer); 
  port ( -- 
    size : in  std_logic_vector(31 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendOutput;
architecture sendOutput_arch of sendOutput is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal size_buffer :  std_logic_vector(31 downto 0);
  signal size_update_enable: Boolean;
  -- output port buffer signals
  signal sendOutput_CP_320_start: Boolean;
  signal sendOutput_CP_320_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_ConvTranspose_output_pipe_222_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_222_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_222_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_222_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_225_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_225_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_225_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_225_inst_ack_1 : boolean;
  signal if_stmt_85_branch_req_0 : boolean;
  signal if_stmt_85_branch_ack_1 : boolean;
  signal if_stmt_85_branch_ack_0 : boolean;
  signal type_cast_112_inst_req_0 : boolean;
  signal type_cast_112_inst_ack_0 : boolean;
  signal type_cast_112_inst_req_1 : boolean;
  signal type_cast_112_inst_ack_1 : boolean;
  signal array_obj_ref_141_index_offset_req_0 : boolean;
  signal array_obj_ref_141_index_offset_ack_0 : boolean;
  signal array_obj_ref_141_index_offset_req_1 : boolean;
  signal array_obj_ref_141_index_offset_ack_1 : boolean;
  signal addr_of_142_final_reg_req_0 : boolean;
  signal addr_of_142_final_reg_ack_0 : boolean;
  signal addr_of_142_final_reg_req_1 : boolean;
  signal addr_of_142_final_reg_ack_1 : boolean;
  signal ptr_deref_146_load_0_req_0 : boolean;
  signal ptr_deref_146_load_0_ack_0 : boolean;
  signal ptr_deref_146_load_0_req_1 : boolean;
  signal ptr_deref_146_load_0_ack_1 : boolean;
  signal type_cast_150_inst_req_0 : boolean;
  signal type_cast_150_inst_ack_0 : boolean;
  signal type_cast_150_inst_req_1 : boolean;
  signal type_cast_150_inst_ack_1 : boolean;
  signal type_cast_160_inst_req_0 : boolean;
  signal type_cast_160_inst_ack_0 : boolean;
  signal type_cast_160_inst_req_1 : boolean;
  signal type_cast_160_inst_ack_1 : boolean;
  signal type_cast_170_inst_req_0 : boolean;
  signal type_cast_170_inst_ack_0 : boolean;
  signal type_cast_170_inst_req_1 : boolean;
  signal type_cast_170_inst_ack_1 : boolean;
  signal type_cast_180_inst_req_0 : boolean;
  signal type_cast_180_inst_ack_0 : boolean;
  signal type_cast_180_inst_req_1 : boolean;
  signal type_cast_180_inst_ack_1 : boolean;
  signal type_cast_190_inst_req_0 : boolean;
  signal type_cast_190_inst_ack_0 : boolean;
  signal type_cast_190_inst_req_1 : boolean;
  signal type_cast_190_inst_ack_1 : boolean;
  signal type_cast_200_inst_req_0 : boolean;
  signal type_cast_200_inst_ack_0 : boolean;
  signal type_cast_200_inst_req_1 : boolean;
  signal type_cast_200_inst_ack_1 : boolean;
  signal type_cast_210_inst_req_0 : boolean;
  signal type_cast_210_inst_ack_0 : boolean;
  signal type_cast_210_inst_req_1 : boolean;
  signal type_cast_210_inst_ack_1 : boolean;
  signal type_cast_220_inst_req_0 : boolean;
  signal type_cast_220_inst_ack_0 : boolean;
  signal type_cast_220_inst_req_1 : boolean;
  signal type_cast_220_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_228_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_228_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_228_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_228_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_231_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_231_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_231_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_231_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_234_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_234_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_234_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_234_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_237_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_237_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_237_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_237_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_240_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_240_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_240_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_240_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_243_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_243_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_243_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_243_inst_ack_1 : boolean;
  signal if_stmt_257_branch_req_0 : boolean;
  signal if_stmt_257_branch_ack_1 : boolean;
  signal if_stmt_257_branch_ack_0 : boolean;
  signal phi_stmt_129_req_0 : boolean;
  signal type_cast_135_inst_req_0 : boolean;
  signal type_cast_135_inst_ack_0 : boolean;
  signal type_cast_135_inst_req_1 : boolean;
  signal type_cast_135_inst_ack_1 : boolean;
  signal phi_stmt_129_req_1 : boolean;
  signal phi_stmt_129_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendOutput_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 32) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= size;
  size_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(tag_length + 31 downto 32) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 31 downto 32);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendOutput_CP_320_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendOutput_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_320_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendOutput_CP_320_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_320_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendOutput_CP_320: Block -- control-path 
    signal sendOutput_CP_320_elements: BooleanArray(59 downto 0);
    -- 
  begin -- 
    sendOutput_CP_320_elements(0) <= sendOutput_CP_320_start;
    sendOutput_CP_320_symbol <= sendOutput_CP_320_elements(59);
    -- CP-element group 0:  branch  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (15) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_78/$entry
      -- CP-element group 0: 	 branch_block_stmt_78/branch_block_stmt_78__entry__
      -- CP-element group 0: 	 branch_block_stmt_78/assign_stmt_84__entry__
      -- CP-element group 0: 	 branch_block_stmt_78/assign_stmt_84__exit__
      -- CP-element group 0: 	 branch_block_stmt_78/if_stmt_85__entry__
      -- CP-element group 0: 	 branch_block_stmt_78/assign_stmt_84/$entry
      -- CP-element group 0: 	 branch_block_stmt_78/assign_stmt_84/$exit
      -- CP-element group 0: 	 branch_block_stmt_78/if_stmt_85_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_78/if_stmt_85_eval_test/$entry
      -- CP-element group 0: 	 branch_block_stmt_78/if_stmt_85_eval_test/$exit
      -- CP-element group 0: 	 branch_block_stmt_78/if_stmt_85_eval_test/branch_req
      -- CP-element group 0: 	 branch_block_stmt_78/R_cmp68_86_place
      -- CP-element group 0: 	 branch_block_stmt_78/if_stmt_85_if_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_78/if_stmt_85_else_link/$entry
      -- 
    branch_req_358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(0), ack => if_stmt_85_branch_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	3 
    -- CP-element group 1: 	4 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 branch_block_stmt_78/merge_stmt_91__exit__
      -- CP-element group 1: 	 branch_block_stmt_78/assign_stmt_97_to_assign_stmt_126__entry__
      -- CP-element group 1: 	 branch_block_stmt_78/if_stmt_85_if_link/$exit
      -- CP-element group 1: 	 branch_block_stmt_78/if_stmt_85_if_link/if_choice_transition
      -- CP-element group 1: 	 branch_block_stmt_78/entry_bbx_xnph
      -- CP-element group 1: 	 branch_block_stmt_78/assign_stmt_97_to_assign_stmt_126/$entry
      -- CP-element group 1: 	 branch_block_stmt_78/assign_stmt_97_to_assign_stmt_126/type_cast_112_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_78/assign_stmt_97_to_assign_stmt_126/type_cast_112_update_start_
      -- CP-element group 1: 	 branch_block_stmt_78/assign_stmt_97_to_assign_stmt_126/type_cast_112_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_78/assign_stmt_97_to_assign_stmt_126/type_cast_112_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_78/assign_stmt_97_to_assign_stmt_126/type_cast_112_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_78/assign_stmt_97_to_assign_stmt_126/type_cast_112_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_78/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_78/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 1: 	 branch_block_stmt_78/merge_stmt_91_PhiReqMerge
      -- CP-element group 1: 	 branch_block_stmt_78/merge_stmt_91_PhiAck/$entry
      -- CP-element group 1: 	 branch_block_stmt_78/merge_stmt_91_PhiAck/$exit
      -- CP-element group 1: 	 branch_block_stmt_78/merge_stmt_91_PhiAck/dummy
      -- 
    if_choice_transition_363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_85_branch_ack_1, ack => sendOutput_CP_320_elements(1)); -- 
    rr_380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(1), ack => type_cast_112_inst_req_0); -- 
    cr_385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(1), ack => type_cast_112_inst_req_1); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	59 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_78/if_stmt_85_else_link/$exit
      -- CP-element group 2: 	 branch_block_stmt_78/if_stmt_85_else_link/else_choice_transition
      -- CP-element group 2: 	 branch_block_stmt_78/entry_forx_xend
      -- CP-element group 2: 	 branch_block_stmt_78/entry_forx_xend_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_78/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_85_branch_ack_0, ack => sendOutput_CP_320_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	1 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_78/assign_stmt_97_to_assign_stmt_126/type_cast_112_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_78/assign_stmt_97_to_assign_stmt_126/type_cast_112_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_78/assign_stmt_97_to_assign_stmt_126/type_cast_112_Sample/ra
      -- 
    ra_381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_112_inst_ack_0, ack => sendOutput_CP_320_elements(3)); -- 
    -- CP-element group 4:  transition  place  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	1 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	53 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_78/assign_stmt_97_to_assign_stmt_126__exit__
      -- CP-element group 4: 	 branch_block_stmt_78/bbx_xnph_forx_xbody
      -- CP-element group 4: 	 branch_block_stmt_78/assign_stmt_97_to_assign_stmt_126/$exit
      -- CP-element group 4: 	 branch_block_stmt_78/assign_stmt_97_to_assign_stmt_126/type_cast_112_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_78/assign_stmt_97_to_assign_stmt_126/type_cast_112_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_78/assign_stmt_97_to_assign_stmt_126/type_cast_112_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_78/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_78/bbx_xnph_forx_xbody_PhiReq/phi_stmt_129/$entry
      -- CP-element group 4: 	 branch_block_stmt_78/bbx_xnph_forx_xbody_PhiReq/phi_stmt_129/phi_stmt_129_sources/$entry
      -- 
    ca_386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_112_inst_ack_1, ack => sendOutput_CP_320_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	58 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	50 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_final_index_sum_regn_sample_complete
      -- CP-element group 5: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_final_index_sum_regn_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_final_index_sum_regn_Sample/ack
      -- 
    ack_415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_141_index_offset_ack_0, ack => sendOutput_CP_320_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	58 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (11) 
      -- CP-element group 6: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/addr_of_142_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_root_address_calculated
      -- CP-element group 6: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_offset_calculated
      -- CP-element group 6: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_final_index_sum_regn_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_final_index_sum_regn_Update/ack
      -- CP-element group 6: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_base_plus_offset/$entry
      -- CP-element group 6: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_base_plus_offset/$exit
      -- CP-element group 6: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_base_plus_offset/sum_rename_req
      -- CP-element group 6: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_base_plus_offset/sum_rename_ack
      -- CP-element group 6: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/addr_of_142_request/$entry
      -- CP-element group 6: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/addr_of_142_request/req
      -- 
    ack_420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_141_index_offset_ack_1, ack => sendOutput_CP_320_elements(6)); -- 
    req_429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(6), ack => addr_of_142_final_reg_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/addr_of_142_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/addr_of_142_request/$exit
      -- CP-element group 7: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/addr_of_142_request/ack
      -- 
    ack_430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_142_final_reg_ack_0, ack => sendOutput_CP_320_elements(7)); -- 
    -- CP-element group 8:  join  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	58 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (24) 
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/addr_of_142_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/addr_of_142_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/addr_of_142_complete/ack
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_base_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_word_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_root_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_base_address_resized
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_base_addr_resize/$entry
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_base_addr_resize/$exit
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_base_addr_resize/base_resize_req
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_base_addr_resize/base_resize_ack
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_base_plus_offset/$entry
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_base_plus_offset/$exit
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_base_plus_offset/sum_rename_req
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_base_plus_offset/sum_rename_ack
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_word_addrgen/$entry
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_word_addrgen/$exit
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_word_addrgen/root_register_req
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_word_addrgen/root_register_ack
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_Sample/word_access_start/$entry
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_Sample/word_access_start/word_0/$entry
      -- CP-element group 8: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_Sample/word_access_start/word_0/rr
      -- 
    ack_435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_142_final_reg_ack_1, ack => sendOutput_CP_320_elements(8)); -- 
    rr_468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(8), ack => ptr_deref_146_load_0_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_Sample/word_access_start/word_0/ra
      -- 
    ra_469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_146_load_0_ack_0, ack => sendOutput_CP_320_elements(9)); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	58 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	17 
    -- CP-element group 10: 	19 
    -- CP-element group 10: 	21 
    -- CP-element group 10: 	23 
    -- CP-element group 10: 	25 
    -- CP-element group 10:  members (33) 
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_Update/ptr_deref_146_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_Update/ptr_deref_146_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_Update/ptr_deref_146_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_Update/ptr_deref_146_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_150_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_150_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_150_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_160_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_160_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_160_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_170_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_170_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_170_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_180_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_180_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_180_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_190_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_190_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_190_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_200_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_200_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_200_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_210_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_210_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_210_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_220_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_220_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_220_Sample/rr
      -- 
    ca_480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_146_load_0_ack_1, ack => sendOutput_CP_320_elements(10)); -- 
    rr_493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(10), ack => type_cast_150_inst_req_0); -- 
    rr_507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(10), ack => type_cast_160_inst_req_0); -- 
    rr_521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(10), ack => type_cast_170_inst_req_0); -- 
    rr_535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(10), ack => type_cast_180_inst_req_0); -- 
    rr_549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(10), ack => type_cast_190_inst_req_0); -- 
    rr_563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(10), ack => type_cast_200_inst_req_0); -- 
    rr_577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(10), ack => type_cast_210_inst_req_0); -- 
    rr_591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(10), ack => type_cast_220_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_150_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_150_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_150_Sample/ra
      -- 
    ra_494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_150_inst_ack_0, ack => sendOutput_CP_320_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	58 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	47 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_150_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_150_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_150_Update/ca
      -- 
    ca_499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_150_inst_ack_1, ack => sendOutput_CP_320_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_160_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_160_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_160_Sample/ra
      -- 
    ra_508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_160_inst_ack_0, ack => sendOutput_CP_320_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	58 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	44 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_160_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_160_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_160_Update/ca
      -- 
    ca_513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_160_inst_ack_1, ack => sendOutput_CP_320_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_170_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_170_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_170_Sample/ra
      -- 
    ra_522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_170_inst_ack_0, ack => sendOutput_CP_320_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	58 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	41 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_170_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_170_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_170_Update/ca
      -- 
    ca_527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_170_inst_ack_1, ack => sendOutput_CP_320_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	10 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_180_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_180_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_180_Sample/ra
      -- 
    ra_536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_180_inst_ack_0, ack => sendOutput_CP_320_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	58 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	38 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_180_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_180_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_180_Update/ca
      -- 
    ca_541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_180_inst_ack_1, ack => sendOutput_CP_320_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	10 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_190_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_190_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_190_Sample/ra
      -- 
    ra_550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_190_inst_ack_0, ack => sendOutput_CP_320_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	58 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	35 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_190_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_190_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_190_Update/ca
      -- 
    ca_555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_190_inst_ack_1, ack => sendOutput_CP_320_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	10 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_200_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_200_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_200_Sample/ra
      -- 
    ra_564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_200_inst_ack_0, ack => sendOutput_CP_320_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	58 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	32 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_200_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_200_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_200_Update/ca
      -- 
    ca_569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_200_inst_ack_1, ack => sendOutput_CP_320_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	10 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_210_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_210_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_210_Sample/ra
      -- 
    ra_578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_210_inst_ack_0, ack => sendOutput_CP_320_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	58 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	29 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_210_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_210_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_210_Update/ca
      -- 
    ca_583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_210_inst_ack_1, ack => sendOutput_CP_320_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	10 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_220_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_220_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_220_Sample/ra
      -- 
    ra_592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_220_inst_ack_0, ack => sendOutput_CP_320_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	58 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_222_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_222_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_222_Sample/req
      -- CP-element group 26: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_220_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_220_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_220_Update/ca
      -- 
    ca_597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_220_inst_ack_1, ack => sendOutput_CP_320_elements(26)); -- 
    req_605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(26), ack => WPIPE_ConvTranspose_output_pipe_222_inst_req_0); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_222_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_222_update_start_
      -- CP-element group 27: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_222_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_222_Sample/ack
      -- CP-element group 27: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_222_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_222_Update/req
      -- 
    ack_606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_222_inst_ack_0, ack => sendOutput_CP_320_elements(27)); -- 
    req_610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(27), ack => WPIPE_ConvTranspose_output_pipe_222_inst_req_1); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_222_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_222_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_222_Update/ack
      -- 
    ack_611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_222_inst_ack_1, ack => sendOutput_CP_320_elements(28)); -- 
    -- CP-element group 29:  join  transition  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	24 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_225_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_225_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_225_Sample/req
      -- 
    req_619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(29), ack => WPIPE_ConvTranspose_output_pipe_225_inst_req_0); -- 
    sendOutput_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_320_elements(24) & sendOutput_CP_320_elements(28);
      gj_sendOutput_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_320_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_225_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_225_update_start_
      -- CP-element group 30: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_225_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_225_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_225_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_225_Update/req
      -- 
    ack_620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_225_inst_ack_0, ack => sendOutput_CP_320_elements(30)); -- 
    req_624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(30), ack => WPIPE_ConvTranspose_output_pipe_225_inst_req_1); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_225_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_225_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_225_Update/ack
      -- 
    ack_625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_225_inst_ack_1, ack => sendOutput_CP_320_elements(31)); -- 
    -- CP-element group 32:  join  transition  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	22 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_228_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_228_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_228_Sample/req
      -- 
    req_633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(32), ack => WPIPE_ConvTranspose_output_pipe_228_inst_req_0); -- 
    sendOutput_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_320_elements(22) & sendOutput_CP_320_elements(31);
      gj_sendOutput_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_320_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_228_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_228_update_start_
      -- CP-element group 33: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_228_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_228_Sample/ack
      -- CP-element group 33: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_228_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_228_Update/req
      -- 
    ack_634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_228_inst_ack_0, ack => sendOutput_CP_320_elements(33)); -- 
    req_638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(33), ack => WPIPE_ConvTranspose_output_pipe_228_inst_req_1); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_228_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_228_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_228_Update/ack
      -- 
    ack_639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_228_inst_ack_1, ack => sendOutput_CP_320_elements(34)); -- 
    -- CP-element group 35:  join  transition  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	20 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_231_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_231_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_231_Sample/req
      -- 
    req_647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(35), ack => WPIPE_ConvTranspose_output_pipe_231_inst_req_0); -- 
    sendOutput_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_320_elements(20) & sendOutput_CP_320_elements(34);
      gj_sendOutput_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_320_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_231_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_231_update_start_
      -- CP-element group 36: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_231_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_231_Sample/ack
      -- CP-element group 36: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_231_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_231_Update/req
      -- 
    ack_648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_231_inst_ack_0, ack => sendOutput_CP_320_elements(36)); -- 
    req_652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(36), ack => WPIPE_ConvTranspose_output_pipe_231_inst_req_1); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_231_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_231_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_231_Update/ack
      -- 
    ack_653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_231_inst_ack_1, ack => sendOutput_CP_320_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	18 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_234_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_234_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_234_Sample/req
      -- 
    req_661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(38), ack => WPIPE_ConvTranspose_output_pipe_234_inst_req_0); -- 
    sendOutput_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_320_elements(18) & sendOutput_CP_320_elements(37);
      gj_sendOutput_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_320_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (6) 
      -- CP-element group 39: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_234_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_234_update_start_
      -- CP-element group 39: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_234_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_234_Sample/ack
      -- CP-element group 39: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_234_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_234_Update/req
      -- 
    ack_662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_234_inst_ack_0, ack => sendOutput_CP_320_elements(39)); -- 
    req_666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(39), ack => WPIPE_ConvTranspose_output_pipe_234_inst_req_1); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_234_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_234_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_234_Update/ack
      -- 
    ack_667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_234_inst_ack_1, ack => sendOutput_CP_320_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	16 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_237_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_237_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_237_Sample/req
      -- 
    req_675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(41), ack => WPIPE_ConvTranspose_output_pipe_237_inst_req_0); -- 
    sendOutput_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_320_elements(16) & sendOutput_CP_320_elements(40);
      gj_sendOutput_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_320_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_237_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_237_update_start_
      -- CP-element group 42: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_237_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_237_Sample/ack
      -- CP-element group 42: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_237_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_237_Update/req
      -- 
    ack_676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_237_inst_ack_0, ack => sendOutput_CP_320_elements(42)); -- 
    req_680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(42), ack => WPIPE_ConvTranspose_output_pipe_237_inst_req_1); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_237_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_237_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_237_Update/ack
      -- 
    ack_681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_237_inst_ack_1, ack => sendOutput_CP_320_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	14 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_240_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_240_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_240_Sample/req
      -- 
    req_689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(44), ack => WPIPE_ConvTranspose_output_pipe_240_inst_req_0); -- 
    sendOutput_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_320_elements(14) & sendOutput_CP_320_elements(43);
      gj_sendOutput_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_320_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_240_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_240_update_start_
      -- CP-element group 45: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_240_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_240_Sample/ack
      -- CP-element group 45: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_240_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_240_Update/req
      -- 
    ack_690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_240_inst_ack_0, ack => sendOutput_CP_320_elements(45)); -- 
    req_694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(45), ack => WPIPE_ConvTranspose_output_pipe_240_inst_req_1); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_240_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_240_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_240_Update/ack
      -- 
    ack_695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_240_inst_ack_1, ack => sendOutput_CP_320_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	12 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_243_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_243_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_243_Sample/req
      -- 
    req_703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(47), ack => WPIPE_ConvTranspose_output_pipe_243_inst_req_0); -- 
    sendOutput_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_320_elements(12) & sendOutput_CP_320_elements(46);
      gj_sendOutput_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_320_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_243_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_243_update_start_
      -- CP-element group 48: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_243_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_243_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_243_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_243_Update/req
      -- 
    ack_704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_243_inst_ack_0, ack => sendOutput_CP_320_elements(48)); -- 
    req_708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(48), ack => WPIPE_ConvTranspose_output_pipe_243_inst_req_1); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_243_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_243_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/WPIPE_ConvTranspose_output_pipe_243_Update/ack
      -- 
    ack_709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_243_inst_ack_1, ack => sendOutput_CP_320_elements(49)); -- 
    -- CP-element group 50:  branch  join  transition  place  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	5 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (10) 
      -- CP-element group 50: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256__exit__
      -- CP-element group 50: 	 branch_block_stmt_78/if_stmt_257__entry__
      -- CP-element group 50: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/$exit
      -- CP-element group 50: 	 branch_block_stmt_78/if_stmt_257_dead_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_78/if_stmt_257_eval_test/$entry
      -- CP-element group 50: 	 branch_block_stmt_78/if_stmt_257_eval_test/$exit
      -- CP-element group 50: 	 branch_block_stmt_78/if_stmt_257_eval_test/branch_req
      -- CP-element group 50: 	 branch_block_stmt_78/R_exitcond1_258_place
      -- CP-element group 50: 	 branch_block_stmt_78/if_stmt_257_if_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_78/if_stmt_257_else_link/$entry
      -- 
    branch_req_717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(50), ack => if_stmt_257_branch_req_0); -- 
    sendOutput_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_320_elements(5) & sendOutput_CP_320_elements(49);
      gj_sendOutput_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_320_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  merge  transition  place  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	59 
    -- CP-element group 51:  members (13) 
      -- CP-element group 51: 	 branch_block_stmt_78/merge_stmt_263__exit__
      -- CP-element group 51: 	 branch_block_stmt_78/forx_xendx_xloopexit_forx_xend
      -- CP-element group 51: 	 branch_block_stmt_78/if_stmt_257_if_link/$exit
      -- CP-element group 51: 	 branch_block_stmt_78/if_stmt_257_if_link/if_choice_transition
      -- CP-element group 51: 	 branch_block_stmt_78/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 51: 	 branch_block_stmt_78/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_78/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 51: 	 branch_block_stmt_78/merge_stmt_263_PhiReqMerge
      -- CP-element group 51: 	 branch_block_stmt_78/merge_stmt_263_PhiAck/$entry
      -- CP-element group 51: 	 branch_block_stmt_78/merge_stmt_263_PhiAck/$exit
      -- CP-element group 51: 	 branch_block_stmt_78/merge_stmt_263_PhiAck/dummy
      -- CP-element group 51: 	 branch_block_stmt_78/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_78/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_257_branch_ack_1, ack => sendOutput_CP_320_elements(51)); -- 
    -- CP-element group 52:  fork  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (12) 
      -- CP-element group 52: 	 branch_block_stmt_78/if_stmt_257_else_link/$exit
      -- CP-element group 52: 	 branch_block_stmt_78/if_stmt_257_else_link/else_choice_transition
      -- CP-element group 52: 	 branch_block_stmt_78/forx_xbody_forx_xbody
      -- CP-element group 52: 	 branch_block_stmt_78/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 52: 	 branch_block_stmt_78/forx_xbody_forx_xbody_PhiReq/phi_stmt_129/$entry
      -- CP-element group 52: 	 branch_block_stmt_78/forx_xbody_forx_xbody_PhiReq/phi_stmt_129/phi_stmt_129_sources/$entry
      -- CP-element group 52: 	 branch_block_stmt_78/forx_xbody_forx_xbody_PhiReq/phi_stmt_129/phi_stmt_129_sources/type_cast_135/$entry
      -- CP-element group 52: 	 branch_block_stmt_78/forx_xbody_forx_xbody_PhiReq/phi_stmt_129/phi_stmt_129_sources/type_cast_135/SplitProtocol/$entry
      -- CP-element group 52: 	 branch_block_stmt_78/forx_xbody_forx_xbody_PhiReq/phi_stmt_129/phi_stmt_129_sources/type_cast_135/SplitProtocol/Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_78/forx_xbody_forx_xbody_PhiReq/phi_stmt_129/phi_stmt_129_sources/type_cast_135/SplitProtocol/Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_78/forx_xbody_forx_xbody_PhiReq/phi_stmt_129/phi_stmt_129_sources/type_cast_135/SplitProtocol/Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_78/forx_xbody_forx_xbody_PhiReq/phi_stmt_129/phi_stmt_129_sources/type_cast_135/SplitProtocol/Update/cr
      -- 
    else_choice_transition_726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_257_branch_ack_0, ack => sendOutput_CP_320_elements(52)); -- 
    rr_770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(52), ack => type_cast_135_inst_req_0); -- 
    cr_775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(52), ack => type_cast_135_inst_req_1); -- 
    -- CP-element group 53:  transition  output  delay-element  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	4 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	57 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_78/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 53: 	 branch_block_stmt_78/bbx_xnph_forx_xbody_PhiReq/phi_stmt_129/$exit
      -- CP-element group 53: 	 branch_block_stmt_78/bbx_xnph_forx_xbody_PhiReq/phi_stmt_129/phi_stmt_129_sources/$exit
      -- CP-element group 53: 	 branch_block_stmt_78/bbx_xnph_forx_xbody_PhiReq/phi_stmt_129/phi_stmt_129_sources/type_cast_133_konst_delay_trans
      -- CP-element group 53: 	 branch_block_stmt_78/bbx_xnph_forx_xbody_PhiReq/phi_stmt_129/phi_stmt_129_req
      -- 
    phi_stmt_129_req_751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_129_req_751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(53), ack => phi_stmt_129_req_0); -- 
    -- Element group sendOutput_CP_320_elements(53) is a control-delay.
    cp_element_53_delay: control_delay_element  generic map(name => " 53_delay", delay_value => 1)  port map(req => sendOutput_CP_320_elements(4), ack => sendOutput_CP_320_elements(53), clk => clk, reset =>reset);
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (2) 
      -- CP-element group 54: 	 branch_block_stmt_78/forx_xbody_forx_xbody_PhiReq/phi_stmt_129/phi_stmt_129_sources/type_cast_135/SplitProtocol/Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_78/forx_xbody_forx_xbody_PhiReq/phi_stmt_129/phi_stmt_129_sources/type_cast_135/SplitProtocol/Sample/ra
      -- 
    ra_771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_135_inst_ack_0, ack => sendOutput_CP_320_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	52 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_78/forx_xbody_forx_xbody_PhiReq/phi_stmt_129/phi_stmt_129_sources/type_cast_135/SplitProtocol/Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_78/forx_xbody_forx_xbody_PhiReq/phi_stmt_129/phi_stmt_129_sources/type_cast_135/SplitProtocol/Update/ca
      -- 
    ca_776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_135_inst_ack_1, ack => sendOutput_CP_320_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (6) 
      -- CP-element group 56: 	 branch_block_stmt_78/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_78/forx_xbody_forx_xbody_PhiReq/phi_stmt_129/$exit
      -- CP-element group 56: 	 branch_block_stmt_78/forx_xbody_forx_xbody_PhiReq/phi_stmt_129/phi_stmt_129_sources/$exit
      -- CP-element group 56: 	 branch_block_stmt_78/forx_xbody_forx_xbody_PhiReq/phi_stmt_129/phi_stmt_129_sources/type_cast_135/$exit
      -- CP-element group 56: 	 branch_block_stmt_78/forx_xbody_forx_xbody_PhiReq/phi_stmt_129/phi_stmt_129_sources/type_cast_135/SplitProtocol/$exit
      -- CP-element group 56: 	 branch_block_stmt_78/forx_xbody_forx_xbody_PhiReq/phi_stmt_129/phi_stmt_129_req
      -- 
    phi_stmt_129_req_777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_129_req_777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(56), ack => phi_stmt_129_req_1); -- 
    sendOutput_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_320_elements(54) & sendOutput_CP_320_elements(55);
      gj_sendOutput_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_320_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  merge  transition  place  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: 	53 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_78/merge_stmt_128_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_78/merge_stmt_128_PhiAck/$entry
      -- 
    sendOutput_CP_320_elements(57) <= OrReduce(sendOutput_CP_320_elements(56) & sendOutput_CP_320_elements(53));
    -- CP-element group 58:  fork  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	5 
    -- CP-element group 58: 	6 
    -- CP-element group 58: 	8 
    -- CP-element group 58: 	10 
    -- CP-element group 58: 	12 
    -- CP-element group 58: 	14 
    -- CP-element group 58: 	16 
    -- CP-element group 58: 	18 
    -- CP-element group 58: 	20 
    -- CP-element group 58: 	22 
    -- CP-element group 58: 	24 
    -- CP-element group 58: 	26 
    -- CP-element group 58:  members (53) 
      -- CP-element group 58: 	 branch_block_stmt_78/merge_stmt_128__exit__
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256__entry__
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/$entry
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/addr_of_142_update_start_
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_final_index_sum_regn_update_start
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_final_index_sum_regn_Sample/req
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_final_index_sum_regn_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/array_obj_ref_141_final_index_sum_regn_Update/req
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/addr_of_142_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/addr_of_142_complete/req
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_update_start_
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_Update/word_access_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_Update/word_access_complete/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/ptr_deref_146_Update/word_access_complete/word_0/cr
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_150_update_start_
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_150_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_150_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_160_update_start_
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_160_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_160_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_170_update_start_
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_170_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_170_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_180_update_start_
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_180_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_180_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_190_update_start_
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_190_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_190_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_200_update_start_
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_200_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_200_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_210_update_start_
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_210_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_210_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_220_update_start_
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_220_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_78/assign_stmt_143_to_assign_stmt_256/type_cast_220_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_78/merge_stmt_128_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_78/merge_stmt_128_PhiAck/phi_stmt_129_ack
      -- 
    phi_stmt_129_ack_782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_129_ack_0, ack => sendOutput_CP_320_elements(58)); -- 
    req_414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(58), ack => array_obj_ref_141_index_offset_req_0); -- 
    req_419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(58), ack => array_obj_ref_141_index_offset_req_1); -- 
    req_434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(58), ack => addr_of_142_final_reg_req_1); -- 
    cr_479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(58), ack => ptr_deref_146_load_0_req_1); -- 
    cr_498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(58), ack => type_cast_150_inst_req_1); -- 
    cr_512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(58), ack => type_cast_160_inst_req_1); -- 
    cr_526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(58), ack => type_cast_170_inst_req_1); -- 
    cr_540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(58), ack => type_cast_180_inst_req_1); -- 
    cr_554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(58), ack => type_cast_190_inst_req_1); -- 
    cr_568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(58), ack => type_cast_200_inst_req_1); -- 
    cr_582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(58), ack => type_cast_210_inst_req_1); -- 
    cr_596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_320_elements(58), ack => type_cast_220_inst_req_1); -- 
    -- CP-element group 59:  merge  transition  place  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	2 
    -- CP-element group 59: 	51 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (16) 
      -- CP-element group 59: 	 $exit
      -- CP-element group 59: 	 branch_block_stmt_78/$exit
      -- CP-element group 59: 	 branch_block_stmt_78/branch_block_stmt_78__exit__
      -- CP-element group 59: 	 branch_block_stmt_78/merge_stmt_265__exit__
      -- CP-element group 59: 	 branch_block_stmt_78/return__
      -- CP-element group 59: 	 branch_block_stmt_78/merge_stmt_267__exit__
      -- CP-element group 59: 	 branch_block_stmt_78/merge_stmt_265_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_78/merge_stmt_265_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_78/merge_stmt_265_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_78/merge_stmt_265_PhiAck/dummy
      -- CP-element group 59: 	 branch_block_stmt_78/return___PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_78/return___PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_78/merge_stmt_267_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_78/merge_stmt_267_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_78/merge_stmt_267_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_78/merge_stmt_267_PhiAck/dummy
      -- 
    sendOutput_CP_320_elements(59) <= OrReduce(sendOutput_CP_320_elements(2) & sendOutput_CP_320_elements(51));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar_140_resized : std_logic_vector(13 downto 0);
    signal R_indvar_140_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_141_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_141_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_141_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_141_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_141_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_141_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_143 : std_logic_vector(31 downto 0);
    signal cmp68_84 : std_logic_vector(0 downto 0);
    signal conv12_161 : std_logic_vector(7 downto 0);
    signal conv18_171 : std_logic_vector(7 downto 0);
    signal conv24_181 : std_logic_vector(7 downto 0);
    signal conv30_191 : std_logic_vector(7 downto 0);
    signal conv36_201 : std_logic_vector(7 downto 0);
    signal conv42_211 : std_logic_vector(7 downto 0);
    signal conv48_221 : std_logic_vector(7 downto 0);
    signal conv_151 : std_logic_vector(7 downto 0);
    signal exitcond1_256 : std_logic_vector(0 downto 0);
    signal iNsTr_1_113 : std_logic_vector(63 downto 0);
    signal indvar_129 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_251 : std_logic_vector(63 downto 0);
    signal ptr_deref_146_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_146_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_146_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_146_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_146_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr15_167 : std_logic_vector(63 downto 0);
    signal shr21_177 : std_logic_vector(63 downto 0);
    signal shr27_187 : std_logic_vector(63 downto 0);
    signal shr33_197 : std_logic_vector(63 downto 0);
    signal shr39_207 : std_logic_vector(63 downto 0);
    signal shr45_217 : std_logic_vector(63 downto 0);
    signal shr9_157 : std_logic_vector(63 downto 0);
    signal shr_97 : std_logic_vector(31 downto 0);
    signal shrx_xop_109 : std_logic_vector(31 downto 0);
    signal tmp4_147 : std_logic_vector(63 downto 0);
    signal tmp72_126 : std_logic_vector(63 downto 0);
    signal tmp_103 : std_logic_vector(0 downto 0);
    signal type_cast_101_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_107_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_117_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_124_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_133_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_135_wire : std_logic_vector(63 downto 0);
    signal type_cast_155_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_165_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_175_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_185_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_195_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_205_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_215_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_249_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_82_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_95_wire_constant : std_logic_vector(31 downto 0);
    signal xx_xop_119 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_141_constant_part_of_offset <= "00000000000000";
    array_obj_ref_141_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_141_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_141_resized_base_address <= "00000000000000";
    ptr_deref_146_word_offset_0 <= "00000000000000";
    type_cast_101_wire_constant <= "00000000000000000000000000000001";
    type_cast_107_wire_constant <= "11111111111111111111111111111111";
    type_cast_117_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_124_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_133_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_155_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_165_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_175_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_185_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_195_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_205_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_215_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_249_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_82_wire_constant <= "00000000000000000000000000000011";
    type_cast_95_wire_constant <= "00000000000000000000000000000010";
    phi_stmt_129: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_133_wire_constant & type_cast_135_wire;
      req <= phi_stmt_129_req_0 & phi_stmt_129_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_129",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_129_ack_0,
          idata => idata,
          odata => indvar_129,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_129
    -- flow-through select operator MUX_125_inst
    tmp72_126 <= xx_xop_119 when (tmp_103(0) /=  '0') else type_cast_124_wire_constant;
    addr_of_142_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_142_final_reg_req_0;
      addr_of_142_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_142_final_reg_req_1;
      addr_of_142_final_reg_ack_1<= rack(0);
      addr_of_142_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_142_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_141_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_143,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_112_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_112_inst_req_0;
      type_cast_112_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_112_inst_req_1;
      type_cast_112_inst_ack_1<= rack(0);
      type_cast_112_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_112_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shrx_xop_109,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_1_113,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_135_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_135_inst_req_0;
      type_cast_135_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_135_inst_req_1;
      type_cast_135_inst_ack_1<= rack(0);
      type_cast_135_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_135_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_251,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_135_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_150_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_150_inst_req_0;
      type_cast_150_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_150_inst_req_1;
      type_cast_150_inst_ack_1<= rack(0);
      type_cast_150_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_150_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp4_147,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_151,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_160_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_160_inst_req_0;
      type_cast_160_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_160_inst_req_1;
      type_cast_160_inst_ack_1<= rack(0);
      type_cast_160_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_160_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr9_157,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_161,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_170_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_170_inst_req_0;
      type_cast_170_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_170_inst_req_1;
      type_cast_170_inst_ack_1<= rack(0);
      type_cast_170_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_170_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr15_167,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv18_171,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_180_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_180_inst_req_0;
      type_cast_180_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_180_inst_req_1;
      type_cast_180_inst_ack_1<= rack(0);
      type_cast_180_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_180_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr21_177,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv24_181,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_190_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_190_inst_req_0;
      type_cast_190_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_190_inst_req_1;
      type_cast_190_inst_ack_1<= rack(0);
      type_cast_190_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_190_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr27_187,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv30_191,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_200_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_200_inst_req_0;
      type_cast_200_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_200_inst_req_1;
      type_cast_200_inst_ack_1<= rack(0);
      type_cast_200_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_200_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr33_197,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv36_201,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_210_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_210_inst_req_0;
      type_cast_210_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_210_inst_req_1;
      type_cast_210_inst_ack_1<= rack(0);
      type_cast_210_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_210_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr39_207,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_211,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_220_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_220_inst_req_0;
      type_cast_220_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_220_inst_req_1;
      type_cast_220_inst_ack_1<= rack(0);
      type_cast_220_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_220_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr45_217,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv48_221,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_141_index_1_rename
    process(R_indvar_140_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_140_resized;
      ov(13 downto 0) := iv;
      R_indvar_140_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_141_index_1_resize
    process(indvar_129) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_129;
      ov := iv(13 downto 0);
      R_indvar_140_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_141_root_address_inst
    process(array_obj_ref_141_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_141_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_141_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_146_addr_0
    process(ptr_deref_146_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_146_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_146_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_146_base_resize
    process(arrayidx_143) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_143;
      ov := iv(13 downto 0);
      ptr_deref_146_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_146_gather_scatter
    process(ptr_deref_146_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_146_data_0;
      ov(63 downto 0) := iv;
      tmp4_147 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_146_root_address_inst
    process(ptr_deref_146_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_146_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_146_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_257_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_256;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_257_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_257_branch_req_0,
          ack0 => if_stmt_257_branch_ack_0,
          ack1 => if_stmt_257_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_85_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp68_84;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_85_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_85_branch_req_0,
          ack0 => if_stmt_85_branch_ack_0,
          ack1 => if_stmt_85_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_108_inst
    process(shr_97) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr_97, type_cast_107_wire_constant, tmp_var);
      shrx_xop_109 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_118_inst
    process(iNsTr_1_113) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_1_113, type_cast_117_wire_constant, tmp_var);
      xx_xop_119 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_250_inst
    process(indvar_129) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_129, type_cast_249_wire_constant, tmp_var);
      indvarx_xnext_251 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_255_inst
    process(indvarx_xnext_251, tmp72_126) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_251, tmp72_126, tmp_var);
      exitcond1_256 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_96_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(size_buffer, type_cast_95_wire_constant, tmp_var);
      shr_97 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_156_inst
    process(tmp4_147) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_147, type_cast_155_wire_constant, tmp_var);
      shr9_157 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_166_inst
    process(tmp4_147) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_147, type_cast_165_wire_constant, tmp_var);
      shr15_167 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_176_inst
    process(tmp4_147) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_147, type_cast_175_wire_constant, tmp_var);
      shr21_177 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_186_inst
    process(tmp4_147) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_147, type_cast_185_wire_constant, tmp_var);
      shr27_187 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_196_inst
    process(tmp4_147) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_147, type_cast_195_wire_constant, tmp_var);
      shr33_197 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_206_inst
    process(tmp4_147) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_147, type_cast_205_wire_constant, tmp_var);
      shr39_207 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_216_inst
    process(tmp4_147) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_147, type_cast_215_wire_constant, tmp_var);
      shr45_217 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_102_inst
    process(shr_97) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_97, type_cast_101_wire_constant, tmp_var);
      tmp_103 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_83_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(size_buffer, type_cast_82_wire_constant, tmp_var);
      cmp68_84 <= tmp_var; --
    end process;
    -- shared split operator group (14) : array_obj_ref_141_index_offset 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_140_scaled;
      array_obj_ref_141_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_141_index_offset_req_0;
      array_obj_ref_141_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_141_index_offset_req_1;
      array_obj_ref_141_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_14_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared load operator group (0) : ptr_deref_146_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_146_load_0_req_0;
      ptr_deref_146_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_146_load_0_req_1;
      ptr_deref_146_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_146_word_address_0;
      ptr_deref_146_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_ConvTranspose_output_pipe_234_inst WPIPE_ConvTranspose_output_pipe_231_inst WPIPE_ConvTranspose_output_pipe_228_inst WPIPE_ConvTranspose_output_pipe_225_inst WPIPE_ConvTranspose_output_pipe_222_inst WPIPE_ConvTranspose_output_pipe_243_inst WPIPE_ConvTranspose_output_pipe_240_inst WPIPE_ConvTranspose_output_pipe_237_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_234_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_231_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_228_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_225_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_222_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_243_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_240_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_237_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_234_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_231_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_228_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_225_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_222_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_243_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_240_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_237_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_234_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_231_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_228_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_225_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_222_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_243_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_240_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_237_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_234_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_231_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_228_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_225_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_222_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_243_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_240_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_237_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv24_181 & conv30_191 & conv36_201 & conv42_211 & conv48_221 & conv_151 & conv12_161 & conv18_171;
      ConvTranspose_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendOutput_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_281_start: Boolean;
  signal timer_CP_281_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_73_load_0_req_0 : boolean;
  signal LOAD_count_73_load_0_ack_0 : boolean;
  signal LOAD_count_73_load_0_req_1 : boolean;
  signal LOAD_count_73_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_281_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_281_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_281_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_281_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_281: Block -- control-path 
    signal timer_CP_281_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_281_elements(0) <= timer_CP_281_start;
    timer_CP_281_symbol <= timer_CP_281_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_74/$entry
      -- CP-element group 0: 	 assign_stmt_74/LOAD_count_73_sample_start_
      -- CP-element group 0: 	 assign_stmt_74/LOAD_count_73_update_start_
      -- CP-element group 0: 	 assign_stmt_74/LOAD_count_73_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_74/LOAD_count_73_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_74/LOAD_count_73_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_74/LOAD_count_73_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_74/LOAD_count_73_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_74/LOAD_count_73_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_74/LOAD_count_73_Update/$entry
      -- CP-element group 0: 	 assign_stmt_74/LOAD_count_73_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_74/LOAD_count_73_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_74/LOAD_count_73_Update/word_access_complete/word_0/cr
      -- 
    cr_313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_281_elements(0), ack => LOAD_count_73_load_0_req_1); -- 
    rr_302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_281_elements(0), ack => LOAD_count_73_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_74/LOAD_count_73_sample_completed_
      -- CP-element group 1: 	 assign_stmt_74/LOAD_count_73_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_74/LOAD_count_73_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_74/LOAD_count_73_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_74/LOAD_count_73_Sample/word_access_start/word_0/ra
      -- 
    ra_303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_73_load_0_ack_0, ack => timer_CP_281_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_74/$exit
      -- CP-element group 2: 	 assign_stmt_74/LOAD_count_73_update_completed_
      -- CP-element group 2: 	 assign_stmt_74/LOAD_count_73_Update/$exit
      -- CP-element group 2: 	 assign_stmt_74/LOAD_count_73_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_74/LOAD_count_73_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_74/LOAD_count_73_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_74/LOAD_count_73_Update/LOAD_count_73_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_74/LOAD_count_73_Update/LOAD_count_73_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_74/LOAD_count_73_Update/LOAD_count_73_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_74/LOAD_count_73_Update/LOAD_count_73_Merge/merge_ack
      -- 
    ca_314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_73_load_0_ack_1, ack => timer_CP_281_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_73_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_73_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_73_word_address_0 <= "0";
    -- equivalence LOAD_count_73_gather_scatter
    process(LOAD_count_73_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_73_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_73_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_73_load_0_req_0;
      LOAD_count_73_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_73_load_0_req_1;
      LOAD_count_73_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_73_word_address_0;
      LOAD_count_73_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(11 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(1 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(1 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      fill_kernel_call_reqs : out  std_logic_vector(0 downto 0);
      fill_kernel_call_acks : in   std_logic_vector(0 downto 0);
      fill_kernel_call_data : out  std_logic_vector(63 downto 0);
      fill_kernel_call_tag  :  out  std_logic_vector(0 downto 0);
      fill_kernel_return_reqs : out  std_logic_vector(0 downto 0);
      fill_kernel_return_acks : in   std_logic_vector(0 downto 0);
      fill_kernel_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_call_acks : in   std_logic_vector(0 downto 0);
      sendOutput_call_data : out  std_logic_vector(31 downto 0);
      sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
      sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_return_acks : in   std_logic_vector(0 downto 0);
      sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module fill_kernel
  component fill_kernel is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(63 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(11 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module fill_kernel
  signal fill_kernel_addr :  std_logic_vector(63 downto 0);
  signal fill_kernel_in_args    : std_logic_vector(63 downto 0);
  signal fill_kernel_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal fill_kernel_tag_out   : std_logic_vector(1 downto 0);
  signal fill_kernel_start_req : std_logic;
  signal fill_kernel_start_ack : std_logic;
  signal fill_kernel_fin_req   : std_logic;
  signal fill_kernel_fin_ack : std_logic;
  -- caller side aggregated signals for module fill_kernel
  signal fill_kernel_call_reqs: std_logic_vector(0 downto 0);
  signal fill_kernel_call_acks: std_logic_vector(0 downto 0);
  signal fill_kernel_return_reqs: std_logic_vector(0 downto 0);
  signal fill_kernel_return_acks: std_logic_vector(0 downto 0);
  signal fill_kernel_call_data: std_logic_vector(63 downto 0);
  signal fill_kernel_call_tag: std_logic_vector(0 downto 0);
  signal fill_kernel_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sendOutput
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendOutput
  signal sendOutput_size :  std_logic_vector(31 downto 0);
  signal sendOutput_in_args    : std_logic_vector(31 downto 0);
  signal sendOutput_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendOutput_tag_out   : std_logic_vector(1 downto 0);
  signal sendOutput_start_req : std_logic;
  signal sendOutput_start_ack : std_logic;
  signal sendOutput_fin_req   : std_logic;
  signal sendOutput_fin_ack : std_logic;
  -- caller side aggregated signals for module sendOutput
  signal sendOutput_call_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_call_acks: std_logic_vector(0 downto 0);
  signal sendOutput_return_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_return_acks: std_logic_vector(0 downto 0);
  signal sendOutput_call_data: std_logic_vector(31 downto 0);
  signal sendOutput_call_tag: std_logic_vector(0 downto 0);
  signal sendOutput_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(1 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(17 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(17 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(13 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(63 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(18 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(1 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      fill_kernel_call_reqs => fill_kernel_call_reqs(0 downto 0),
      fill_kernel_call_acks => fill_kernel_call_acks(0 downto 0),
      fill_kernel_call_data => fill_kernel_call_data(63 downto 0),
      fill_kernel_call_tag => fill_kernel_call_tag(0 downto 0),
      fill_kernel_return_reqs => fill_kernel_return_reqs(0 downto 0),
      fill_kernel_return_acks => fill_kernel_return_acks(0 downto 0),
      fill_kernel_return_tag => fill_kernel_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      sendOutput_call_reqs => sendOutput_call_reqs(0 downto 0),
      sendOutput_call_acks => sendOutput_call_acks(0 downto 0),
      sendOutput_call_data => sendOutput_call_data(31 downto 0),
      sendOutput_call_tag => sendOutput_call_tag(0 downto 0),
      sendOutput_return_reqs => sendOutput_return_reqs(0 downto 0),
      sendOutput_return_acks => sendOutput_return_acks(0 downto 0),
      sendOutput_return_tag => sendOutput_return_tag(0 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module fill_kernel
  fill_kernel_addr <= fill_kernel_in_args(63 downto 0);
  -- call arbiter for module fill_kernel
  fill_kernel_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => fill_kernel_call_reqs,
      call_acks => fill_kernel_call_acks,
      return_reqs => fill_kernel_return_reqs,
      return_acks => fill_kernel_return_acks,
      call_data  => fill_kernel_call_data,
      call_tag  => fill_kernel_call_tag,
      return_tag  => fill_kernel_return_tag,
      call_mtag => fill_kernel_tag_in,
      return_mtag => fill_kernel_tag_out,
      call_mreq => fill_kernel_start_req,
      call_mack => fill_kernel_start_ack,
      return_mreq => fill_kernel_fin_req,
      return_mack => fill_kernel_fin_ack,
      call_mdata => fill_kernel_in_args,
      clk => clk, 
      reset => reset --
    ); --
  fill_kernel_instance:fill_kernel-- 
    generic map(tag_length => 2)
    port map(-- 
      addr => fill_kernel_addr,
      start_req => fill_kernel_start_req,
      start_ack => fill_kernel_start_ack,
      fin_req => fill_kernel_fin_req,
      fin_ack => fill_kernel_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(11 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(0 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(1 downto 1),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(1 downto 1),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(15 downto 8),
      tag_in => fill_kernel_tag_in,
      tag_out => fill_kernel_tag_out-- 
    ); -- 
  -- module sendOutput
  sendOutput_size <= sendOutput_in_args(31 downto 0);
  -- call arbiter for module sendOutput
  sendOutput_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendOutput_call_reqs,
      call_acks => sendOutput_call_acks,
      return_reqs => sendOutput_return_reqs,
      return_acks => sendOutput_return_acks,
      call_data  => sendOutput_call_data,
      call_tag  => sendOutput_call_tag,
      return_tag  => sendOutput_return_tag,
      call_mtag => sendOutput_tag_in,
      return_mtag => sendOutput_tag_out,
      call_mreq => sendOutput_start_req,
      call_mack => sendOutput_start_ack,
      return_mreq => sendOutput_fin_req,
      return_mack => sendOutput_fin_ack,
      call_mdata => sendOutput_in_args,
      clk => clk, 
      reset => reset --
    ); --
  sendOutput_instance:sendOutput-- 
    generic map(tag_length => 2)
    port map(-- 
      size => sendOutput_size,
      start_req => sendOutput_start_req,
      start_ack => sendOutput_start_ack,
      fin_req => sendOutput_fin_req,
      fin_ack => sendOutput_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(18 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(1 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      tag_in => sendOutput_tag_in,
      tag_out => sendOutput_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(0 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(0 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 2,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  dummyROM_memory_space_0: dummy_read_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_2: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_stores => 1,
      addr_width => 12,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
