-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_34_start: Boolean;
  signal convTranspose_CP_34_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal WPIPE_Block2_start_1081_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_746_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_746_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_746_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1031_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_539_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_746_inst_req_0 : boolean;
  signal addr_of_694_final_reg_req_0 : boolean;
  signal WPIPE_Block1_start_1063_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_593_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_593_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1075_inst_req_1 : boolean;
  signal WPIPE_Block0_start_978_inst_req_1 : boolean;
  signal if_stmt_637_branch_req_0 : boolean;
  signal WPIPE_Block2_start_1084_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1056_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1034_inst_req_1 : boolean;
  signal type_cast_615_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1002_inst_ack_0 : boolean;
  signal type_cast_615_inst_req_1 : boolean;
  signal type_cast_597_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_593_inst_ack_0 : boolean;
  signal type_cast_543_inst_ack_1 : boolean;
  signal type_cast_597_inst_req_0 : boolean;
  signal type_cast_543_inst_req_1 : boolean;
  signal type_cast_543_inst_ack_0 : boolean;
  signal type_cast_543_inst_req_0 : boolean;
  signal array_obj_ref_693_index_offset_req_1 : boolean;
  signal type_cast_1417_inst_ack_0 : boolean;
  signal ptr_deref_623_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_40_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_40_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_40_inst_req_1 : boolean;
  signal ptr_deref_623_store_0_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_40_inst_ack_1 : boolean;
  signal type_cast_714_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_593_inst_req_0 : boolean;
  signal type_cast_44_inst_req_0 : boolean;
  signal type_cast_44_inst_ack_0 : boolean;
  signal type_cast_44_inst_req_1 : boolean;
  signal type_cast_44_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1087_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1013_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_993_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_140_inst_ack_1 : boolean;
  signal type_cast_144_inst_req_0 : boolean;
  signal WPIPE_Block0_start_978_inst_ack_1 : boolean;
  signal type_cast_144_inst_ack_0 : boolean;
  signal type_cast_714_inst_req_0 : boolean;
  signal type_cast_57_inst_req_0 : boolean;
  signal type_cast_57_inst_ack_0 : boolean;
  signal type_cast_57_inst_req_1 : boolean;
  signal type_cast_57_inst_ack_1 : boolean;
  signal type_cast_664_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_65_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_65_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_697_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_65_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_65_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_728_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1084_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_993_inst_req_0 : boolean;
  signal type_cast_615_inst_ack_0 : boolean;
  signal array_obj_ref_693_index_offset_ack_0 : boolean;
  signal type_cast_69_inst_req_0 : boolean;
  signal type_cast_69_inst_ack_0 : boolean;
  signal type_cast_69_inst_req_1 : boolean;
  signal type_cast_69_inst_ack_1 : boolean;
  signal type_cast_664_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_697_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_78_inst_req_0 : boolean;
  signal ptr_deref_623_store_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_78_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_78_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_78_inst_ack_1 : boolean;
  signal type_cast_1417_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_710_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_710_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1063_inst_ack_0 : boolean;
  signal type_cast_615_inst_req_0 : boolean;
  signal array_obj_ref_693_index_offset_req_0 : boolean;
  signal type_cast_82_inst_req_0 : boolean;
  signal ptr_deref_623_store_0_req_0 : boolean;
  signal type_cast_82_inst_ack_0 : boolean;
  signal type_cast_82_inst_req_1 : boolean;
  signal type_cast_82_inst_ack_1 : boolean;
  signal type_cast_664_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_90_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_90_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_90_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_90_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_728_inst_req_1 : boolean;
  signal type_cast_94_inst_req_0 : boolean;
  signal type_cast_94_inst_ack_0 : boolean;
  signal type_cast_94_inst_req_1 : boolean;
  signal type_cast_94_inst_ack_1 : boolean;
  signal type_cast_714_inst_ack_1 : boolean;
  signal type_cast_732_inst_ack_1 : boolean;
  signal type_cast_664_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_103_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_103_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_103_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1056_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_103_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_710_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_710_inst_req_0 : boolean;
  signal WPIPE_Block0_start_993_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1075_inst_ack_1 : boolean;
  signal type_cast_107_inst_req_0 : boolean;
  signal type_cast_107_inst_ack_0 : boolean;
  signal type_cast_107_inst_req_1 : boolean;
  signal type_cast_107_inst_ack_1 : boolean;
  signal type_cast_714_inst_req_1 : boolean;
  signal WPIPE_Block0_start_978_inst_ack_0 : boolean;
  signal type_cast_732_inst_req_1 : boolean;
  signal type_cast_579_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1016_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1302_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_697_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_115_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_115_inst_ack_0 : boolean;
  signal type_cast_579_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_115_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_115_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_993_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1016_inst_req_0 : boolean;
  signal type_cast_119_inst_req_0 : boolean;
  signal type_cast_119_inst_ack_0 : boolean;
  signal type_cast_119_inst_req_1 : boolean;
  signal type_cast_119_inst_ack_1 : boolean;
  signal addr_of_694_final_reg_ack_1 : boolean;
  signal WPIPE_Block2_start_1090_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_697_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1069_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1019_inst_req_0 : boolean;
  signal type_cast_132_inst_req_0 : boolean;
  signal type_cast_132_inst_ack_0 : boolean;
  signal type_cast_132_inst_req_1 : boolean;
  signal type_cast_132_inst_ack_1 : boolean;
  signal addr_of_694_final_reg_req_1 : boolean;
  signal WPIPE_Block1_start_1069_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_140_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_140_inst_ack_0 : boolean;
  signal type_cast_579_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_140_inst_req_1 : boolean;
  signal type_cast_345_inst_req_1 : boolean;
  signal type_cast_345_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1022_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_354_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_354_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_354_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_354_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1022_inst_ack_1 : boolean;
  signal type_cast_1387_inst_ack_1 : boolean;
  signal type_cast_144_inst_req_1 : boolean;
  signal type_cast_144_inst_ack_1 : boolean;
  signal type_cast_732_inst_ack_0 : boolean;
  signal type_cast_579_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_153_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_153_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_153_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_153_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1090_inst_req_0 : boolean;
  signal WPIPE_Block0_start_978_inst_req_0 : boolean;
  signal type_cast_157_inst_req_0 : boolean;
  signal type_cast_157_inst_ack_0 : boolean;
  signal type_cast_157_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1002_inst_req_0 : boolean;
  signal type_cast_157_inst_ack_1 : boolean;
  signal type_cast_732_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_165_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_165_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_165_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_165_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_728_inst_ack_0 : boolean;
  signal type_cast_169_inst_req_0 : boolean;
  signal type_cast_169_inst_ack_0 : boolean;
  signal type_cast_169_inst_req_1 : boolean;
  signal type_cast_169_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1066_inst_ack_1 : boolean;
  signal addr_of_694_final_reg_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_178_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_178_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_178_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_178_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_539_inst_ack_0 : boolean;
  signal type_cast_182_inst_req_0 : boolean;
  signal type_cast_182_inst_ack_0 : boolean;
  signal type_cast_182_inst_req_1 : boolean;
  signal type_cast_182_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_575_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_190_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_190_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_575_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_190_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_190_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_728_inst_req_0 : boolean;
  signal type_cast_701_inst_ack_1 : boolean;
  signal type_cast_701_inst_req_1 : boolean;
  signal WPIPE_Block0_start_987_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1019_inst_ack_0 : boolean;
  signal type_cast_194_inst_req_0 : boolean;
  signal type_cast_194_inst_ack_0 : boolean;
  signal type_cast_194_inst_req_1 : boolean;
  signal ptr_deref_1373_load_0_ack_1 : boolean;
  signal type_cast_194_inst_ack_1 : boolean;
  signal if_stmt_637_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_203_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_203_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_575_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_203_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_203_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_984_inst_ack_1 : boolean;
  signal type_cast_207_inst_req_0 : boolean;
  signal type_cast_207_inst_ack_0 : boolean;
  signal type_cast_207_inst_req_1 : boolean;
  signal type_cast_207_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_575_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_611_inst_ack_1 : boolean;
  signal type_cast_216_inst_req_0 : boolean;
  signal type_cast_216_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_539_inst_req_0 : boolean;
  signal type_cast_216_inst_req_1 : boolean;
  signal WPIPE_Block0_start_987_inst_ack_0 : boolean;
  signal type_cast_216_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1019_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_611_inst_req_1 : boolean;
  signal type_cast_220_inst_req_0 : boolean;
  signal type_cast_220_inst_ack_0 : boolean;
  signal type_cast_220_inst_req_1 : boolean;
  signal type_cast_220_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1019_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_611_inst_ack_0 : boolean;
  signal type_cast_224_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1056_inst_req_1 : boolean;
  signal type_cast_224_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1016_inst_ack_0 : boolean;
  signal type_cast_224_inst_req_1 : boolean;
  signal type_cast_224_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1063_inst_req_1 : boolean;
  signal type_cast_561_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_611_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1063_inst_ack_1 : boolean;
  signal type_cast_261_inst_req_0 : boolean;
  signal type_cast_261_inst_ack_0 : boolean;
  signal type_cast_261_inst_req_1 : boolean;
  signal type_cast_261_inst_ack_1 : boolean;
  signal type_cast_561_inst_req_1 : boolean;
  signal type_cast_265_inst_req_0 : boolean;
  signal type_cast_265_inst_ack_0 : boolean;
  signal type_cast_265_inst_req_1 : boolean;
  signal type_cast_265_inst_ack_1 : boolean;
  signal type_cast_561_inst_ack_0 : boolean;
  signal type_cast_269_inst_req_0 : boolean;
  signal type_cast_269_inst_ack_0 : boolean;
  signal type_cast_269_inst_req_1 : boolean;
  signal type_cast_269_inst_ack_1 : boolean;
  signal type_cast_561_inst_req_0 : boolean;
  signal type_cast_273_inst_req_0 : boolean;
  signal type_cast_273_inst_ack_0 : boolean;
  signal type_cast_273_inst_req_1 : boolean;
  signal type_cast_273_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_987_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_291_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_291_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_291_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1056_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_291_inst_ack_1 : boolean;
  signal type_cast_701_inst_ack_0 : boolean;
  signal type_cast_701_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1034_inst_req_0 : boolean;
  signal type_cast_295_inst_req_0 : boolean;
  signal type_cast_295_inst_ack_0 : boolean;
  signal type_cast_295_inst_req_1 : boolean;
  signal type_cast_295_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_557_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_304_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_304_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_557_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_304_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_304_inst_ack_1 : boolean;
  signal type_cast_597_inst_ack_1 : boolean;
  signal type_cast_308_inst_req_0 : boolean;
  signal type_cast_308_inst_ack_0 : boolean;
  signal type_cast_308_inst_req_1 : boolean;
  signal type_cast_308_inst_ack_1 : boolean;
  signal if_stmt_637_branch_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_557_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_ack_1 : boolean;
  signal type_cast_597_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1034_inst_ack_0 : boolean;
  signal type_cast_320_inst_req_0 : boolean;
  signal ptr_deref_1373_load_0_req_1 : boolean;
  signal type_cast_320_inst_ack_0 : boolean;
  signal type_cast_320_inst_req_1 : boolean;
  signal type_cast_320_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_557_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_329_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_329_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_329_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_329_inst_ack_1 : boolean;
  signal array_obj_ref_693_index_offset_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_539_inst_ack_1 : boolean;
  signal type_cast_333_inst_req_0 : boolean;
  signal type_cast_333_inst_ack_0 : boolean;
  signal type_cast_333_inst_req_1 : boolean;
  signal type_cast_333_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1034_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_341_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_341_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_341_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_341_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1022_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1022_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_987_inst_ack_1 : boolean;
  signal type_cast_345_inst_req_0 : boolean;
  signal type_cast_345_inst_ack_0 : boolean;
  signal type_cast_358_inst_req_0 : boolean;
  signal type_cast_358_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_981_inst_req_0 : boolean;
  signal type_cast_358_inst_req_1 : boolean;
  signal type_cast_358_inst_ack_1 : boolean;
  signal type_cast_1417_inst_req_0 : boolean;
  signal WPIPE_Block0_start_996_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_ack_0 : boolean;
  signal type_cast_1417_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1302_inst_req_0 : boolean;
  signal type_cast_370_inst_req_0 : boolean;
  signal type_cast_370_inst_ack_0 : boolean;
  signal type_cast_370_inst_req_1 : boolean;
  signal type_cast_370_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_996_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_379_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_379_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_379_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_379_inst_ack_1 : boolean;
  signal type_cast_383_inst_req_0 : boolean;
  signal type_cast_383_inst_ack_0 : boolean;
  signal type_cast_383_inst_req_1 : boolean;
  signal type_cast_383_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1002_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_391_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_391_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_996_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_391_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_391_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_996_inst_ack_1 : boolean;
  signal type_cast_395_inst_req_0 : boolean;
  signal type_cast_395_inst_ack_0 : boolean;
  signal type_cast_395_inst_req_1 : boolean;
  signal type_cast_395_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_404_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_404_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1025_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_404_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_404_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1299_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1025_inst_ack_0 : boolean;
  signal type_cast_408_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1025_inst_req_1 : boolean;
  signal type_cast_408_inst_ack_0 : boolean;
  signal type_cast_408_inst_req_1 : boolean;
  signal type_cast_408_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_981_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1025_inst_ack_1 : boolean;
  signal if_stmt_421_branch_req_0 : boolean;
  signal if_stmt_421_branch_ack_1 : boolean;
  signal if_stmt_421_branch_ack_0 : boolean;
  signal if_stmt_436_branch_req_0 : boolean;
  signal if_stmt_436_branch_ack_1 : boolean;
  signal if_stmt_436_branch_ack_0 : boolean;
  signal type_cast_457_inst_req_0 : boolean;
  signal type_cast_457_inst_ack_0 : boolean;
  signal type_cast_457_inst_req_1 : boolean;
  signal type_cast_457_inst_ack_1 : boolean;
  signal array_obj_ref_486_index_offset_req_0 : boolean;
  signal array_obj_ref_486_index_offset_ack_0 : boolean;
  signal array_obj_ref_486_index_offset_req_1 : boolean;
  signal array_obj_ref_486_index_offset_ack_1 : boolean;
  signal addr_of_487_final_reg_req_0 : boolean;
  signal addr_of_487_final_reg_ack_0 : boolean;
  signal addr_of_487_final_reg_req_1 : boolean;
  signal addr_of_487_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_490_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_490_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_490_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_490_inst_ack_1 : boolean;
  signal type_cast_494_inst_req_0 : boolean;
  signal type_cast_494_inst_ack_0 : boolean;
  signal type_cast_494_inst_req_1 : boolean;
  signal type_cast_494_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1016_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_503_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_503_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_503_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_503_inst_ack_1 : boolean;
  signal type_cast_507_inst_req_0 : boolean;
  signal type_cast_507_inst_ack_0 : boolean;
  signal type_cast_507_inst_req_1 : boolean;
  signal type_cast_507_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_521_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_521_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_521_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_521_inst_ack_1 : boolean;
  signal type_cast_525_inst_req_0 : boolean;
  signal type_cast_525_inst_ack_0 : boolean;
  signal type_cast_525_inst_req_1 : boolean;
  signal type_cast_525_inst_ack_1 : boolean;
  signal type_cast_750_inst_req_0 : boolean;
  signal type_cast_750_inst_ack_0 : boolean;
  signal type_cast_750_inst_req_1 : boolean;
  signal type_cast_750_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1087_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1066_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_764_inst_req_0 : boolean;
  signal type_cast_1054_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_764_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1081_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_764_inst_req_1 : boolean;
  signal type_cast_1054_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_764_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1458_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1084_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1084_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1287_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1013_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1072_inst_ack_1 : boolean;
  signal type_cast_768_inst_req_0 : boolean;
  signal type_cast_768_inst_ack_0 : boolean;
  signal type_cast_768_inst_req_1 : boolean;
  signal type_cast_768_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_990_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1066_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_782_inst_req_0 : boolean;
  signal type_cast_1054_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_782_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_990_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_782_inst_req_1 : boolean;
  signal type_cast_1054_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_782_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1075_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1013_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1072_inst_req_1 : boolean;
  signal type_cast_786_inst_req_0 : boolean;
  signal type_cast_786_inst_ack_0 : boolean;
  signal type_cast_786_inst_req_1 : boolean;
  signal type_cast_786_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1066_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_800_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_800_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1081_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_800_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_800_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1075_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1013_inst_req_0 : boolean;
  signal type_cast_804_inst_req_0 : boolean;
  signal type_cast_804_inst_ack_0 : boolean;
  signal type_cast_804_inst_req_1 : boolean;
  signal type_cast_804_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1078_inst_ack_1 : boolean;
  signal type_cast_1387_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1290_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_818_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1043_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_818_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_990_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1081_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_818_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1043_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_818_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1458_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1290_inst_ack_0 : boolean;
  signal type_cast_822_inst_req_0 : boolean;
  signal type_cast_822_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1072_inst_ack_0 : boolean;
  signal type_cast_822_inst_req_1 : boolean;
  signal type_cast_822_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1087_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1078_inst_req_1 : boolean;
  signal type_cast_1061_inst_ack_1 : boolean;
  signal type_cast_1061_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1043_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1043_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1031_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1072_inst_req_0 : boolean;
  signal ptr_deref_830_store_0_req_0 : boolean;
  signal WPIPE_Block0_start_1010_inst_ack_1 : boolean;
  signal ptr_deref_830_store_0_ack_0 : boolean;
  signal WPIPE_Block0_start_984_inst_req_1 : boolean;
  signal WPIPE_Block0_start_999_inst_ack_1 : boolean;
  signal ptr_deref_830_store_0_req_1 : boolean;
  signal WPIPE_Block0_start_1010_inst_req_1 : boolean;
  signal ptr_deref_830_store_0_ack_1 : boolean;
  signal if_stmt_844_branch_req_0 : boolean;
  signal WPIPE_Block0_start_1010_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1031_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_984_inst_ack_0 : boolean;
  signal if_stmt_844_branch_ack_1 : boolean;
  signal WPIPE_Block1_start_1031_inst_req_0 : boolean;
  signal WPIPE_Block0_start_984_inst_req_0 : boolean;
  signal if_stmt_844_branch_ack_0 : boolean;
  signal WPIPE_Block0_start_999_inst_req_1 : boolean;
  signal type_cast_855_inst_req_0 : boolean;
  signal type_cast_855_inst_ack_0 : boolean;
  signal type_cast_855_inst_req_1 : boolean;
  signal type_cast_855_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1087_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1078_inst_ack_0 : boolean;
  signal type_cast_1339_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1010_inst_req_0 : boolean;
  signal type_cast_859_inst_req_0 : boolean;
  signal type_cast_859_inst_ack_0 : boolean;
  signal type_cast_859_inst_req_1 : boolean;
  signal type_cast_859_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1078_inst_req_0 : boolean;
  signal type_cast_1061_inst_ack_0 : boolean;
  signal type_cast_1061_inst_req_0 : boolean;
  signal type_cast_863_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1040_inst_ack_1 : boolean;
  signal type_cast_863_inst_ack_0 : boolean;
  signal type_cast_863_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1040_inst_req_1 : boolean;
  signal type_cast_863_inst_ack_1 : boolean;
  signal if_stmt_881_branch_req_0 : boolean;
  signal if_stmt_881_branch_ack_1 : boolean;
  signal if_stmt_881_branch_ack_0 : boolean;
  signal WPIPE_Block1_start_1028_inst_ack_1 : boolean;
  signal type_cast_908_inst_req_0 : boolean;
  signal type_cast_908_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1028_inst_req_1 : boolean;
  signal type_cast_908_inst_req_1 : boolean;
  signal type_cast_908_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1090_inst_ack_1 : boolean;
  signal type_cast_1339_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1287_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1006_inst_ack_1 : boolean;
  signal array_obj_ref_937_index_offset_req_0 : boolean;
  signal WPIPE_Block1_start_1040_inst_ack_0 : boolean;
  signal array_obj_ref_937_index_offset_ack_0 : boolean;
  signal WPIPE_Block0_start_990_inst_req_0 : boolean;
  signal array_obj_ref_937_index_offset_req_1 : boolean;
  signal WPIPE_Block1_start_1040_inst_req_0 : boolean;
  signal array_obj_ref_937_index_offset_ack_1 : boolean;
  signal WPIPE_Block0_start_1006_inst_req_1 : boolean;
  signal addr_of_938_final_reg_req_0 : boolean;
  signal addr_of_938_final_reg_ack_0 : boolean;
  signal addr_of_938_final_reg_req_1 : boolean;
  signal addr_of_938_final_reg_ack_1 : boolean;
  signal WPIPE_Block2_start_1090_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1299_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1302_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1006_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1028_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1037_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1037_inst_req_1 : boolean;
  signal WPIPE_Block0_start_999_inst_ack_0 : boolean;
  signal ptr_deref_941_store_0_req_0 : boolean;
  signal WPIPE_Block0_start_1006_inst_req_0 : boolean;
  signal ptr_deref_941_store_0_ack_0 : boolean;
  signal WPIPE_Block1_start_1028_inst_req_0 : boolean;
  signal WPIPE_Block0_start_999_inst_req_0 : boolean;
  signal ptr_deref_941_store_0_req_1 : boolean;
  signal ptr_deref_941_store_0_ack_1 : boolean;
  signal WPIPE_Block0_start_981_inst_ack_1 : boolean;
  signal if_stmt_956_branch_req_0 : boolean;
  signal WPIPE_Block0_start_981_inst_req_1 : boolean;
  signal if_stmt_956_branch_ack_1 : boolean;
  signal if_stmt_956_branch_ack_0 : boolean;
  signal call_stmt_967_call_req_0 : boolean;
  signal call_stmt_967_call_ack_0 : boolean;
  signal WPIPE_Block1_start_1069_inst_ack_1 : boolean;
  signal call_stmt_967_call_req_1 : boolean;
  signal call_stmt_967_call_ack_1 : boolean;
  signal type_cast_1397_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1037_inst_ack_0 : boolean;
  signal type_cast_972_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1037_inst_req_0 : boolean;
  signal type_cast_972_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1069_inst_req_1 : boolean;
  signal type_cast_972_inst_req_1 : boolean;
  signal type_cast_972_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1002_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_975_inst_req_0 : boolean;
  signal WPIPE_Block0_start_975_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_975_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1302_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_975_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1093_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1093_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1093_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1093_inst_ack_1 : boolean;
  signal type_cast_1387_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1455_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1096_inst_req_0 : boolean;
  signal ptr_deref_1373_load_0_ack_0 : boolean;
  signal WPIPE_Block2_start_1096_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1455_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1096_inst_req_1 : boolean;
  signal ptr_deref_1373_load_0_req_0 : boolean;
  signal WPIPE_Block2_start_1096_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1452_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1452_inst_req_1 : boolean;
  signal type_cast_1339_inst_ack_0 : boolean;
  signal type_cast_1387_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1099_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1099_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1299_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1099_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1099_inst_ack_1 : boolean;
  signal type_cast_1339_inst_req_0 : boolean;
  signal type_cast_1427_inst_ack_1 : boolean;
  signal type_cast_1110_inst_req_0 : boolean;
  signal type_cast_1110_inst_ack_0 : boolean;
  signal type_cast_1427_inst_req_1 : boolean;
  signal type_cast_1110_inst_req_1 : boolean;
  signal type_cast_1110_inst_ack_1 : boolean;
  signal type_cast_1407_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1112_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1112_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1299_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1112_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1112_inst_ack_1 : boolean;
  signal type_cast_1117_inst_req_0 : boolean;
  signal type_cast_1117_inst_ack_0 : boolean;
  signal type_cast_1117_inst_req_1 : boolean;
  signal type_cast_1117_inst_ack_1 : boolean;
  signal type_cast_1377_inst_ack_1 : boolean;
  signal type_cast_1377_inst_req_1 : boolean;
  signal type_cast_1407_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1455_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1119_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1119_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1119_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1119_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1452_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1452_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1122_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1122_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1455_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1122_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1122_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1458_inst_ack_0 : boolean;
  signal type_cast_1427_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1125_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1125_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1125_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1125_inst_ack_1 : boolean;
  signal type_cast_1377_inst_ack_0 : boolean;
  signal type_cast_1407_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1128_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1128_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1128_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1128_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1458_inst_req_0 : boolean;
  signal type_cast_1377_inst_req_0 : boolean;
  signal type_cast_1407_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1131_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1131_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1296_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1131_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1131_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1134_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1134_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1296_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1134_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1134_inst_ack_1 : boolean;
  signal if_stmt_1312_branch_ack_0 : boolean;
  signal WPIPE_Block3_start_1137_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1137_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1137_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1137_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1140_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1140_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1140_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1140_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1449_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1449_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1143_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1143_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1296_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1143_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1143_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1296_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1449_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1449_inst_req_0 : boolean;
  signal if_stmt_1312_branch_ack_1 : boolean;
  signal WPIPE_Block3_start_1146_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1146_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1146_inst_req_1 : boolean;
  signal addr_of_1369_final_reg_ack_1 : boolean;
  signal WPIPE_Block3_start_1146_inst_ack_1 : boolean;
  signal type_cast_1427_inst_req_0 : boolean;
  signal if_stmt_1312_branch_req_0 : boolean;
  signal WPIPE_Block3_start_1149_inst_req_0 : boolean;
  signal addr_of_1369_final_reg_req_1 : boolean;
  signal WPIPE_Block3_start_1149_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1149_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1149_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1152_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1152_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1152_inst_req_1 : boolean;
  signal addr_of_1369_final_reg_ack_0 : boolean;
  signal WPIPE_Block3_start_1152_inst_ack_1 : boolean;
  signal type_cast_1447_inst_ack_1 : boolean;
  signal type_cast_1447_inst_req_1 : boolean;
  signal type_cast_1397_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1155_inst_req_0 : boolean;
  signal addr_of_1369_final_reg_req_0 : boolean;
  signal WPIPE_Block3_start_1155_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1155_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1155_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1293_inst_ack_1 : boolean;
  signal type_cast_1447_inst_ack_0 : boolean;
  signal type_cast_1447_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1308_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1308_inst_req_1 : boolean;
  signal type_cast_1166_inst_req_0 : boolean;
  signal type_cast_1166_inst_ack_0 : boolean;
  signal type_cast_1166_inst_req_1 : boolean;
  signal type_cast_1166_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1293_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1308_inst_ack_0 : boolean;
  signal type_cast_1397_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1168_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1168_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1168_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1168_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1293_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1308_inst_req_0 : boolean;
  signal type_cast_1173_inst_req_0 : boolean;
  signal type_cast_1173_inst_ack_0 : boolean;
  signal type_cast_1173_inst_req_1 : boolean;
  signal array_obj_ref_1368_index_offset_ack_1 : boolean;
  signal type_cast_1173_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1293_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1175_inst_req_0 : boolean;
  signal array_obj_ref_1368_index_offset_req_1 : boolean;
  signal WPIPE_Block3_start_1175_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1175_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1175_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1305_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1305_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1178_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1178_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1178_inst_req_1 : boolean;
  signal array_obj_ref_1368_index_offset_ack_0 : boolean;
  signal WPIPE_Block3_start_1178_inst_ack_1 : boolean;
  signal type_cast_1437_inst_ack_1 : boolean;
  signal type_cast_1437_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1305_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1181_inst_req_0 : boolean;
  signal array_obj_ref_1368_index_offset_req_0 : boolean;
  signal WPIPE_Block3_start_1181_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1181_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1181_inst_ack_1 : boolean;
  signal type_cast_1437_inst_ack_0 : boolean;
  signal type_cast_1437_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1305_inst_req_0 : boolean;
  signal type_cast_1397_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1184_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1184_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1290_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1184_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1184_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1290_inst_req_1 : boolean;
  signal RPIPE_Block0_done_1189_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1189_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_1189_inst_req_1 : boolean;
  signal RPIPE_Block0_done_1189_inst_ack_1 : boolean;
  signal RPIPE_Block1_done_1192_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1192_inst_ack_0 : boolean;
  signal RPIPE_Block1_done_1192_inst_req_1 : boolean;
  signal RPIPE_Block1_done_1192_inst_ack_1 : boolean;
  signal RPIPE_Block2_done_1195_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1195_inst_ack_0 : boolean;
  signal RPIPE_Block2_done_1195_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1195_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1198_inst_req_0 : boolean;
  signal RPIPE_Block3_done_1198_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1198_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1198_inst_ack_1 : boolean;
  signal call_stmt_1202_call_req_0 : boolean;
  signal call_stmt_1202_call_ack_0 : boolean;
  signal call_stmt_1202_call_req_1 : boolean;
  signal call_stmt_1202_call_ack_1 : boolean;
  signal type_cast_1206_inst_req_0 : boolean;
  signal type_cast_1206_inst_ack_0 : boolean;
  signal type_cast_1206_inst_req_1 : boolean;
  signal type_cast_1206_inst_ack_1 : boolean;
  signal type_cast_1215_inst_req_0 : boolean;
  signal type_cast_1215_inst_ack_0 : boolean;
  signal type_cast_1215_inst_req_1 : boolean;
  signal type_cast_1215_inst_ack_1 : boolean;
  signal type_cast_1225_inst_req_0 : boolean;
  signal type_cast_1225_inst_ack_0 : boolean;
  signal type_cast_1225_inst_req_1 : boolean;
  signal type_cast_1225_inst_ack_1 : boolean;
  signal type_cast_1235_inst_req_0 : boolean;
  signal type_cast_1235_inst_ack_0 : boolean;
  signal type_cast_1235_inst_req_1 : boolean;
  signal type_cast_1235_inst_ack_1 : boolean;
  signal type_cast_1245_inst_req_0 : boolean;
  signal type_cast_1245_inst_ack_0 : boolean;
  signal type_cast_1245_inst_req_1 : boolean;
  signal type_cast_1245_inst_ack_1 : boolean;
  signal type_cast_1255_inst_req_0 : boolean;
  signal type_cast_1255_inst_ack_0 : boolean;
  signal type_cast_1255_inst_req_1 : boolean;
  signal type_cast_1255_inst_ack_1 : boolean;
  signal type_cast_1265_inst_req_0 : boolean;
  signal type_cast_1265_inst_ack_0 : boolean;
  signal type_cast_1265_inst_req_1 : boolean;
  signal type_cast_1265_inst_ack_1 : boolean;
  signal type_cast_1275_inst_req_0 : boolean;
  signal type_cast_1275_inst_ack_0 : boolean;
  signal type_cast_1275_inst_req_1 : boolean;
  signal type_cast_1275_inst_ack_1 : boolean;
  signal type_cast_1285_inst_req_0 : boolean;
  signal type_cast_1285_inst_ack_0 : boolean;
  signal type_cast_1285_inst_req_1 : boolean;
  signal type_cast_1285_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1287_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1287_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1461_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1461_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1461_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1461_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1464_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1464_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1464_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1464_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1467_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1467_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1467_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1467_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1470_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1470_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1470_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1470_inst_ack_1 : boolean;
  signal if_stmt_1484_branch_req_0 : boolean;
  signal if_stmt_1484_branch_ack_1 : boolean;
  signal if_stmt_1484_branch_ack_0 : boolean;
  signal phi_stmt_474_req_0 : boolean;
  signal type_cast_480_inst_req_0 : boolean;
  signal type_cast_480_inst_ack_0 : boolean;
  signal type_cast_480_inst_req_1 : boolean;
  signal type_cast_480_inst_ack_1 : boolean;
  signal phi_stmt_474_req_1 : boolean;
  signal phi_stmt_474_ack_0 : boolean;
  signal phi_stmt_681_req_0 : boolean;
  signal type_cast_687_inst_req_0 : boolean;
  signal type_cast_687_inst_ack_0 : boolean;
  signal type_cast_687_inst_req_1 : boolean;
  signal type_cast_687_inst_ack_1 : boolean;
  signal phi_stmt_681_req_1 : boolean;
  signal phi_stmt_681_ack_0 : boolean;
  signal phi_stmt_925_req_1 : boolean;
  signal type_cast_928_inst_req_0 : boolean;
  signal type_cast_928_inst_ack_0 : boolean;
  signal type_cast_928_inst_req_1 : boolean;
  signal type_cast_928_inst_ack_1 : boolean;
  signal phi_stmt_925_req_0 : boolean;
  signal phi_stmt_925_ack_0 : boolean;
  signal phi_stmt_1356_req_0 : boolean;
  signal type_cast_1362_inst_req_0 : boolean;
  signal type_cast_1362_inst_ack_0 : boolean;
  signal type_cast_1362_inst_req_1 : boolean;
  signal type_cast_1362_inst_ack_1 : boolean;
  signal phi_stmt_1356_req_1 : boolean;
  signal phi_stmt_1356_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_34_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_34_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_34_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_34_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_34: Block -- control-path 
    signal convTranspose_CP_34_elements: BooleanArray(497 downto 0);
    -- 
  begin -- 
    convTranspose_CP_34_elements(0) <= convTranspose_CP_34_start;
    convTranspose_CP_34_symbol <= convTranspose_CP_34_elements(497);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	59 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	68 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	62 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	71 
    -- CP-element group 0: 	74 
    -- CP-element group 0: 	77 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	85 
    -- CP-element group 0: 	89 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	101 
    -- CP-element group 0: 	105 
    -- CP-element group 0: 	109 
    -- CP-element group 0: 	113 
    -- CP-element group 0: 	117 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0:  members (101) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_38/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/branch_block_stmt_38__entry__
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420__entry__
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Update/cr
      -- 
    rr_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => RPIPE_ConvTranspose_input_pipe_40_inst_req_0); -- 
    cr_151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_44_inst_req_1); -- 
    cr_179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_57_inst_req_1); -- 
    cr_207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_69_inst_req_1); -- 
    cr_235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_82_inst_req_1); -- 
    cr_263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_94_inst_req_1); -- 
    cr_291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_107_inst_req_1); -- 
    cr_319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_119_inst_req_1); -- 
    cr_347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_132_inst_req_1); -- 
    cr_753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_345_inst_req_1); -- 
    cr_375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_144_inst_req_1); -- 
    cr_403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_157_inst_req_1); -- 
    cr_431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_169_inst_req_1); -- 
    cr_459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_182_inst_req_1); -- 
    cr_487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_194_inst_req_1); -- 
    cr_515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_207_inst_req_1); -- 
    cr_529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_216_inst_req_1); -- 
    cr_543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_220_inst_req_1); -- 
    cr_557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_224_inst_req_1); -- 
    cr_571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_261_inst_req_1); -- 
    cr_585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_265_inst_req_1); -- 
    cr_599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_269_inst_req_1); -- 
    cr_613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_273_inst_req_1); -- 
    cr_641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_295_inst_req_1); -- 
    cr_669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_308_inst_req_1); -- 
    cr_697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_320_inst_req_1); -- 
    cr_725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_333_inst_req_1); -- 
    cr_781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_358_inst_req_1); -- 
    cr_809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_370_inst_req_1); -- 
    cr_837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_383_inst_req_1); -- 
    cr_865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_395_inst_req_1); -- 
    cr_893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_408_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_update_start_
      -- CP-element group 1: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Update/cr
      -- 
    ra_133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_40_inst_ack_0, ack => convTranspose_CP_34_elements(1)); -- 
    cr_137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(1), ack => RPIPE_ConvTranspose_input_pipe_40_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_sample_start_
      -- 
    ca_138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_40_inst_ack_1, ack => convTranspose_CP_34_elements(2)); -- 
    rr_146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(2), ack => type_cast_44_inst_req_0); -- 
    rr_160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(2), ack => RPIPE_ConvTranspose_input_pipe_53_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Sample/ra
      -- 
    ra_147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_44_inst_ack_0, ack => convTranspose_CP_34_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	57 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Update/ca
      -- 
    ca_152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_44_inst_ack_1, ack => convTranspose_CP_34_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Update/cr
      -- CP-element group 5: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_update_start_
      -- 
    ra_161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_53_inst_ack_0, ack => convTranspose_CP_34_elements(5)); -- 
    cr_165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(5), ack => RPIPE_ConvTranspose_input_pipe_53_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Sample/rr
      -- 
    ca_166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_53_inst_ack_1, ack => convTranspose_CP_34_elements(6)); -- 
    rr_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(6), ack => type_cast_57_inst_req_0); -- 
    rr_188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(6), ack => RPIPE_ConvTranspose_input_pipe_65_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Sample/ra
      -- 
    ra_175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_57_inst_ack_0, ack => convTranspose_CP_34_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	57 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Update/ca
      -- 
    ca_180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_57_inst_ack_1, ack => convTranspose_CP_34_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_update_start_
      -- CP-element group 9: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Update/cr
      -- 
    ra_189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_65_inst_ack_0, ack => convTranspose_CP_34_elements(9)); -- 
    cr_193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(9), ack => RPIPE_ConvTranspose_input_pipe_65_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Sample/rr
      -- 
    ca_194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_65_inst_ack_1, ack => convTranspose_CP_34_elements(10)); -- 
    rr_202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(10), ack => type_cast_69_inst_req_0); -- 
    rr_216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(10), ack => RPIPE_ConvTranspose_input_pipe_78_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Sample/ra
      -- 
    ra_203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_69_inst_ack_0, ack => convTranspose_CP_34_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	60 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Update/ca
      -- 
    ca_208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_69_inst_ack_1, ack => convTranspose_CP_34_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_update_start_
      -- CP-element group 13: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Update/cr
      -- 
    ra_217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_78_inst_ack_0, ack => convTranspose_CP_34_elements(13)); -- 
    cr_221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(13), ack => RPIPE_ConvTranspose_input_pipe_78_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Sample/rr
      -- 
    ca_222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_78_inst_ack_1, ack => convTranspose_CP_34_elements(14)); -- 
    rr_230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(14), ack => type_cast_82_inst_req_0); -- 
    rr_244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(14), ack => RPIPE_ConvTranspose_input_pipe_90_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Sample/ra
      -- 
    ra_231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_82_inst_ack_0, ack => convTranspose_CP_34_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	60 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Update/ca
      -- 
    ca_236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_82_inst_ack_1, ack => convTranspose_CP_34_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_update_start_
      -- CP-element group 17: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Update/cr
      -- 
    ra_245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_90_inst_ack_0, ack => convTranspose_CP_34_elements(17)); -- 
    cr_249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(17), ack => RPIPE_ConvTranspose_input_pipe_90_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Sample/rr
      -- 
    ca_250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_90_inst_ack_1, ack => convTranspose_CP_34_elements(18)); -- 
    rr_258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(18), ack => type_cast_94_inst_req_0); -- 
    rr_272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(18), ack => RPIPE_ConvTranspose_input_pipe_103_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Sample/ra
      -- 
    ra_259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_94_inst_ack_0, ack => convTranspose_CP_34_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	63 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Update/ca
      -- 
    ca_264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_94_inst_ack_1, ack => convTranspose_CP_34_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_update_start_
      -- CP-element group 21: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Update/cr
      -- 
    ra_273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_103_inst_ack_0, ack => convTranspose_CP_34_elements(21)); -- 
    cr_277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(21), ack => RPIPE_ConvTranspose_input_pipe_103_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Sample/rr
      -- 
    ca_278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_103_inst_ack_1, ack => convTranspose_CP_34_elements(22)); -- 
    rr_286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(22), ack => type_cast_107_inst_req_0); -- 
    rr_300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(22), ack => RPIPE_ConvTranspose_input_pipe_115_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Sample/ra
      -- 
    ra_287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_107_inst_ack_0, ack => convTranspose_CP_34_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	63 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Update/ca
      -- 
    ca_292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_107_inst_ack_1, ack => convTranspose_CP_34_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_update_start_
      -- CP-element group 25: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Update/cr
      -- 
    ra_301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_115_inst_ack_0, ack => convTranspose_CP_34_elements(25)); -- 
    cr_305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(25), ack => RPIPE_ConvTranspose_input_pipe_115_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Sample/rr
      -- 
    ca_306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_115_inst_ack_1, ack => convTranspose_CP_34_elements(26)); -- 
    rr_314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(26), ack => type_cast_119_inst_req_0); -- 
    rr_328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(26), ack => RPIPE_ConvTranspose_input_pipe_128_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Sample/ra
      -- 
    ra_315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_119_inst_ack_0, ack => convTranspose_CP_34_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	66 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Update/ca
      -- 
    ca_320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_119_inst_ack_1, ack => convTranspose_CP_34_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_update_start_
      -- CP-element group 29: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Update/cr
      -- 
    ra_329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_128_inst_ack_0, ack => convTranspose_CP_34_elements(29)); -- 
    cr_333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(29), ack => RPIPE_ConvTranspose_input_pipe_128_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Sample/rr
      -- 
    ca_334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_128_inst_ack_1, ack => convTranspose_CP_34_elements(30)); -- 
    rr_342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(30), ack => type_cast_132_inst_req_0); -- 
    rr_356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(30), ack => RPIPE_ConvTranspose_input_pipe_140_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Sample/ra
      -- 
    ra_343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_132_inst_ack_0, ack => convTranspose_CP_34_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	66 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Update/ca
      -- 
    ca_348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_132_inst_ack_1, ack => convTranspose_CP_34_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_update_start_
      -- CP-element group 33: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Update/cr
      -- 
    ra_357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_140_inst_ack_0, ack => convTranspose_CP_34_elements(33)); -- 
    cr_361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(33), ack => RPIPE_ConvTranspose_input_pipe_140_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Sample/rr
      -- 
    ca_362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_140_inst_ack_1, ack => convTranspose_CP_34_elements(34)); -- 
    rr_370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(34), ack => type_cast_144_inst_req_0); -- 
    rr_384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(34), ack => RPIPE_ConvTranspose_input_pipe_153_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Sample/ra
      -- 
    ra_371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_144_inst_ack_0, ack => convTranspose_CP_34_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	69 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Update/ca
      -- 
    ca_376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_144_inst_ack_1, ack => convTranspose_CP_34_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_update_start_
      -- CP-element group 37: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Update/cr
      -- 
    ra_385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_153_inst_ack_0, ack => convTranspose_CP_34_elements(37)); -- 
    cr_389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(37), ack => RPIPE_ConvTranspose_input_pipe_153_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Sample/rr
      -- 
    ca_390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_153_inst_ack_1, ack => convTranspose_CP_34_elements(38)); -- 
    rr_398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(38), ack => type_cast_157_inst_req_0); -- 
    rr_412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(38), ack => RPIPE_ConvTranspose_input_pipe_165_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Sample/ra
      -- 
    ra_399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_157_inst_ack_0, ack => convTranspose_CP_34_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	69 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Update/ca
      -- 
    ca_404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_157_inst_ack_1, ack => convTranspose_CP_34_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_update_start_
      -- CP-element group 41: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Update/cr
      -- 
    ra_413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_165_inst_ack_0, ack => convTranspose_CP_34_elements(41)); -- 
    cr_417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(41), ack => RPIPE_ConvTranspose_input_pipe_165_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	45 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Sample/rr
      -- 
    ca_418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_165_inst_ack_1, ack => convTranspose_CP_34_elements(42)); -- 
    rr_426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(42), ack => type_cast_169_inst_req_0); -- 
    rr_440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(42), ack => RPIPE_ConvTranspose_input_pipe_178_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Sample/ra
      -- 
    ra_427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_169_inst_ack_0, ack => convTranspose_CP_34_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	72 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Update/ca
      -- 
    ca_432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_169_inst_ack_1, ack => convTranspose_CP_34_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_update_start_
      -- CP-element group 45: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Update/cr
      -- 
    ra_441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_178_inst_ack_0, ack => convTranspose_CP_34_elements(45)); -- 
    cr_445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(45), ack => RPIPE_ConvTranspose_input_pipe_178_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	49 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Sample/rr
      -- 
    ca_446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_178_inst_ack_1, ack => convTranspose_CP_34_elements(46)); -- 
    rr_454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(46), ack => type_cast_182_inst_req_0); -- 
    rr_468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(46), ack => RPIPE_ConvTranspose_input_pipe_190_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Sample/ra
      -- 
    ra_455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_182_inst_ack_0, ack => convTranspose_CP_34_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	72 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Update/ca
      -- 
    ca_460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_182_inst_ack_1, ack => convTranspose_CP_34_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_update_start_
      -- CP-element group 49: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Update/cr
      -- 
    ra_469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_190_inst_ack_0, ack => convTranspose_CP_34_elements(49)); -- 
    cr_473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(49), ack => RPIPE_ConvTranspose_input_pipe_190_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Sample/rr
      -- 
    ca_474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_190_inst_ack_1, ack => convTranspose_CP_34_elements(50)); -- 
    rr_496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(50), ack => RPIPE_ConvTranspose_input_pipe_203_inst_req_0); -- 
    rr_482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(50), ack => type_cast_194_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Sample/ra
      -- 
    ra_483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_194_inst_ack_0, ack => convTranspose_CP_34_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	75 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Update/ca
      -- 
    ca_488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_194_inst_ack_1, ack => convTranspose_CP_34_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_update_start_
      -- CP-element group 53: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Update/cr
      -- 
    ra_497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_203_inst_ack_0, ack => convTranspose_CP_34_elements(53)); -- 
    cr_501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(53), ack => RPIPE_ConvTranspose_input_pipe_203_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	78 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Sample/rr
      -- 
    ca_502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_203_inst_ack_1, ack => convTranspose_CP_34_elements(54)); -- 
    rr_510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(54), ack => type_cast_207_inst_req_0); -- 
    rr_622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(54), ack => RPIPE_ConvTranspose_input_pipe_291_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Sample/ra
      -- 
    ra_511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_207_inst_ack_0, ack => convTranspose_CP_34_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	75 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Update/ca
      -- 
    ca_516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_207_inst_ack_1, ack => convTranspose_CP_34_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	4 
    -- CP-element group 57: 	8 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Sample/rr
      -- 
    rr_524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(57), ack => type_cast_216_inst_req_0); -- 
    convTranspose_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(4) & convTranspose_CP_34_elements(8);
      gj_convTranspose_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Sample/ra
      -- 
    ra_525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_216_inst_ack_0, ack => convTranspose_CP_34_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	0 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	118 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Update/ca
      -- 
    ca_530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_216_inst_ack_1, ack => convTranspose_CP_34_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	12 
    -- CP-element group 60: 	16 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Sample/rr
      -- 
    rr_538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(60), ack => type_cast_220_inst_req_0); -- 
    convTranspose_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(12) & convTranspose_CP_34_elements(16);
      gj_convTranspose_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Sample/ra
      -- 
    ra_539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_220_inst_ack_0, ack => convTranspose_CP_34_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	0 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	118 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Update/ca
      -- 
    ca_544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_220_inst_ack_1, ack => convTranspose_CP_34_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	20 
    -- CP-element group 63: 	24 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Sample/rr
      -- 
    rr_552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(63), ack => type_cast_224_inst_req_0); -- 
    convTranspose_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(20) & convTranspose_CP_34_elements(24);
      gj_convTranspose_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Sample/ra
      -- 
    ra_553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_224_inst_ack_0, ack => convTranspose_CP_34_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	118 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Update/ca
      -- 
    ca_558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_224_inst_ack_1, ack => convTranspose_CP_34_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	28 
    -- CP-element group 66: 	32 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Sample/rr
      -- 
    rr_566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(66), ack => type_cast_261_inst_req_0); -- 
    convTranspose_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(28) & convTranspose_CP_34_elements(32);
      gj_convTranspose_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Sample/ra
      -- 
    ra_567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_261_inst_ack_0, ack => convTranspose_CP_34_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	0 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	118 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Update/ca
      -- 
    ca_572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_261_inst_ack_1, ack => convTranspose_CP_34_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	40 
    -- CP-element group 69: 	36 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Sample/rr
      -- 
    rr_580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(69), ack => type_cast_265_inst_req_0); -- 
    convTranspose_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(40) & convTranspose_CP_34_elements(36);
      gj_convTranspose_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Sample/ra
      -- 
    ra_581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_265_inst_ack_0, ack => convTranspose_CP_34_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	0 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	118 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Update/ca
      -- 
    ca_586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_265_inst_ack_1, ack => convTranspose_CP_34_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	48 
    -- CP-element group 72: 	44 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Sample/rr
      -- 
    rr_594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(72), ack => type_cast_269_inst_req_0); -- 
    convTranspose_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(48) & convTranspose_CP_34_elements(44);
      gj_convTranspose_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Sample/ra
      -- 
    ra_595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_269_inst_ack_0, ack => convTranspose_CP_34_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	0 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	118 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Update/ca
      -- 
    ca_600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_269_inst_ack_1, ack => convTranspose_CP_34_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	56 
    -- CP-element group 75: 	52 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Sample/rr
      -- 
    rr_608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(75), ack => type_cast_273_inst_req_0); -- 
    convTranspose_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(56) & convTranspose_CP_34_elements(52);
      gj_convTranspose_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Sample/ra
      -- 
    ra_609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_273_inst_ack_0, ack => convTranspose_CP_34_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	0 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	118 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Update/ca
      -- 
    ca_614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_273_inst_ack_1, ack => convTranspose_CP_34_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	54 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_update_start_
      -- CP-element group 78: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Update/cr
      -- 
    ra_623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_291_inst_ack_0, ack => convTranspose_CP_34_elements(78)); -- 
    cr_627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(78), ack => RPIPE_ConvTranspose_input_pipe_291_inst_req_1); -- 
    -- CP-element group 79:  fork  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	82 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Sample/rr
      -- 
    ca_628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_291_inst_ack_1, ack => convTranspose_CP_34_elements(79)); -- 
    rr_636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(79), ack => type_cast_295_inst_req_0); -- 
    rr_650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(79), ack => RPIPE_ConvTranspose_input_pipe_304_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Sample/ra
      -- 
    ra_637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_295_inst_ack_0, ack => convTranspose_CP_34_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	118 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Update/ca
      -- 
    ca_642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_295_inst_ack_1, ack => convTranspose_CP_34_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_update_start_
      -- CP-element group 82: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Update/cr
      -- 
    ra_651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_304_inst_ack_0, ack => convTranspose_CP_34_elements(82)); -- 
    cr_655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(82), ack => RPIPE_ConvTranspose_input_pipe_304_inst_req_1); -- 
    -- CP-element group 83:  fork  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	86 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Sample/rr
      -- 
    ca_656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_304_inst_ack_1, ack => convTranspose_CP_34_elements(83)); -- 
    rr_664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(83), ack => type_cast_308_inst_req_0); -- 
    rr_678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(83), ack => RPIPE_ConvTranspose_input_pipe_316_inst_req_0); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Sample/ra
      -- 
    ra_665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_308_inst_ack_0, ack => convTranspose_CP_34_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	0 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	118 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Update/ca
      -- 
    ca_670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_308_inst_ack_1, ack => convTranspose_CP_34_elements(85)); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	83 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_update_start_
      -- CP-element group 86: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Update/cr
      -- 
    ra_679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_316_inst_ack_0, ack => convTranspose_CP_34_elements(86)); -- 
    cr_683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(86), ack => RPIPE_ConvTranspose_input_pipe_316_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Sample/rr
      -- 
    ca_684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_316_inst_ack_1, ack => convTranspose_CP_34_elements(87)); -- 
    rr_692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(87), ack => type_cast_320_inst_req_0); -- 
    rr_706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(87), ack => RPIPE_ConvTranspose_input_pipe_329_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Sample/ra
      -- 
    ra_693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_320_inst_ack_0, ack => convTranspose_CP_34_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	0 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	118 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Update/ca
      -- 
    ca_698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_320_inst_ack_1, ack => convTranspose_CP_34_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_update_start_
      -- CP-element group 90: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Update/cr
      -- 
    ra_707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_329_inst_ack_0, ack => convTranspose_CP_34_elements(90)); -- 
    cr_711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(90), ack => RPIPE_ConvTranspose_input_pipe_329_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Sample/rr
      -- 
    ca_712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_329_inst_ack_1, ack => convTranspose_CP_34_elements(91)); -- 
    rr_720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(91), ack => type_cast_333_inst_req_0); -- 
    rr_734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(91), ack => RPIPE_ConvTranspose_input_pipe_341_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Sample/ra
      -- 
    ra_721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_333_inst_ack_0, ack => convTranspose_CP_34_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	118 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Update/ca
      -- 
    ca_726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_333_inst_ack_1, ack => convTranspose_CP_34_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_update_start_
      -- CP-element group 94: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Update/cr
      -- 
    ra_735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_341_inst_ack_0, ack => convTranspose_CP_34_elements(94)); -- 
    cr_739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(94), ack => RPIPE_ConvTranspose_input_pipe_341_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Sample/rr
      -- 
    ca_740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_341_inst_ack_1, ack => convTranspose_CP_34_elements(95)); -- 
    rr_748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(95), ack => type_cast_345_inst_req_0); -- 
    rr_762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(95), ack => RPIPE_ConvTranspose_input_pipe_354_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Sample/ra
      -- 
    ra_749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_345_inst_ack_0, ack => convTranspose_CP_34_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	118 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_update_completed_
      -- 
    ca_754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_345_inst_ack_1, ack => convTranspose_CP_34_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_update_start_
      -- CP-element group 98: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Update/cr
      -- 
    ra_763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_354_inst_ack_0, ack => convTranspose_CP_34_elements(98)); -- 
    cr_767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(98), ack => RPIPE_ConvTranspose_input_pipe_354_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (9) 
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Sample/rr
      -- 
    ca_768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_354_inst_ack_1, ack => convTranspose_CP_34_elements(99)); -- 
    rr_776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(99), ack => type_cast_358_inst_req_0); -- 
    rr_790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(99), ack => RPIPE_ConvTranspose_input_pipe_366_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Sample/ra
      -- 
    ra_777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_358_inst_ack_0, ack => convTranspose_CP_34_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	0 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	118 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Update/ca
      -- 
    ca_782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_358_inst_ack_1, ack => convTranspose_CP_34_elements(101)); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (6) 
      -- CP-element group 102: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_update_start_
      -- CP-element group 102: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Update/cr
      -- 
    ra_791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_366_inst_ack_0, ack => convTranspose_CP_34_elements(102)); -- 
    cr_795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(102), ack => RPIPE_ConvTranspose_input_pipe_366_inst_req_1); -- 
    -- CP-element group 103:  fork  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: 	106 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Sample/rr
      -- 
    ca_796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_366_inst_ack_1, ack => convTranspose_CP_34_elements(103)); -- 
    rr_804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(103), ack => type_cast_370_inst_req_0); -- 
    rr_818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(103), ack => RPIPE_ConvTranspose_input_pipe_379_inst_req_0); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Sample/ra
      -- 
    ra_805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_370_inst_ack_0, ack => convTranspose_CP_34_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	0 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	118 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Update/ca
      -- 
    ca_810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_370_inst_ack_1, ack => convTranspose_CP_34_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	103 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_update_start_
      -- CP-element group 106: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Update/cr
      -- 
    ra_819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_379_inst_ack_0, ack => convTranspose_CP_34_elements(106)); -- 
    cr_823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(106), ack => RPIPE_ConvTranspose_input_pipe_379_inst_req_1); -- 
    -- CP-element group 107:  fork  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Sample/rr
      -- 
    ca_824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_379_inst_ack_1, ack => convTranspose_CP_34_elements(107)); -- 
    rr_832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(107), ack => type_cast_383_inst_req_0); -- 
    rr_846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(107), ack => RPIPE_ConvTranspose_input_pipe_391_inst_req_0); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Sample/ra
      -- 
    ra_833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_383_inst_ack_0, ack => convTranspose_CP_34_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	0 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	118 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Update/ca
      -- 
    ca_838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_383_inst_ack_1, ack => convTranspose_CP_34_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_update_start_
      -- CP-element group 110: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Update/cr
      -- 
    ra_847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_391_inst_ack_0, ack => convTranspose_CP_34_elements(110)); -- 
    cr_851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(110), ack => RPIPE_ConvTranspose_input_pipe_391_inst_req_1); -- 
    -- CP-element group 111:  fork  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Sample/rr
      -- 
    ca_852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_391_inst_ack_1, ack => convTranspose_CP_34_elements(111)); -- 
    rr_860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(111), ack => type_cast_395_inst_req_0); -- 
    rr_874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(111), ack => RPIPE_ConvTranspose_input_pipe_404_inst_req_0); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Sample/ra
      -- 
    ra_861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_395_inst_ack_0, ack => convTranspose_CP_34_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	0 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	118 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Update/ca
      -- 
    ca_866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_395_inst_ack_1, ack => convTranspose_CP_34_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	111 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_update_start_
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Update/cr
      -- 
    ra_875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_404_inst_ack_0, ack => convTranspose_CP_34_elements(114)); -- 
    cr_879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(114), ack => RPIPE_ConvTranspose_input_pipe_404_inst_req_1); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Sample/rr
      -- 
    ca_880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_404_inst_ack_1, ack => convTranspose_CP_34_elements(115)); -- 
    rr_888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(115), ack => type_cast_408_inst_req_0); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Sample/ra
      -- 
    ra_889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_408_inst_ack_0, ack => convTranspose_CP_34_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	0 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Update/ca
      -- 
    ca_894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_408_inst_ack_1, ack => convTranspose_CP_34_elements(117)); -- 
    -- CP-element group 118:  branch  join  transition  place  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	59 
    -- CP-element group 118: 	65 
    -- CP-element group 118: 	68 
    -- CP-element group 118: 	62 
    -- CP-element group 118: 	71 
    -- CP-element group 118: 	74 
    -- CP-element group 118: 	77 
    -- CP-element group 118: 	81 
    -- CP-element group 118: 	85 
    -- CP-element group 118: 	89 
    -- CP-element group 118: 	93 
    -- CP-element group 118: 	97 
    -- CP-element group 118: 	101 
    -- CP-element group 118: 	105 
    -- CP-element group 118: 	109 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (10) 
      -- CP-element group 118: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420__exit__
      -- CP-element group 118: 	 branch_block_stmt_38/if_stmt_421__entry__
      -- CP-element group 118: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/$exit
      -- CP-element group 118: 	 branch_block_stmt_38/if_stmt_421_dead_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_38/if_stmt_421_eval_test/$entry
      -- CP-element group 118: 	 branch_block_stmt_38/if_stmt_421_eval_test/$exit
      -- CP-element group 118: 	 branch_block_stmt_38/if_stmt_421_eval_test/branch_req
      -- CP-element group 118: 	 branch_block_stmt_38/R_cmp513_422_place
      -- CP-element group 118: 	 branch_block_stmt_38/if_stmt_421_if_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_38/if_stmt_421_else_link/$entry
      -- 
    branch_req_902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(118), ack => if_stmt_421_branch_req_0); -- 
    convTranspose_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(59) & convTranspose_CP_34_elements(65) & convTranspose_CP_34_elements(68) & convTranspose_CP_34_elements(62) & convTranspose_CP_34_elements(71) & convTranspose_CP_34_elements(74) & convTranspose_CP_34_elements(77) & convTranspose_CP_34_elements(81) & convTranspose_CP_34_elements(85) & convTranspose_CP_34_elements(89) & convTranspose_CP_34_elements(93) & convTranspose_CP_34_elements(97) & convTranspose_CP_34_elements(101) & convTranspose_CP_34_elements(105) & convTranspose_CP_34_elements(109) & convTranspose_CP_34_elements(113) & convTranspose_CP_34_elements(117);
      gj_convTranspose_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	123 
    -- CP-element group 119: 	124 
    -- CP-element group 119:  members (18) 
      -- CP-element group 119: 	 branch_block_stmt_38/merge_stmt_442__exit__
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471__entry__
      -- CP-element group 119: 	 branch_block_stmt_38/if_stmt_421_if_link/$exit
      -- CP-element group 119: 	 branch_block_stmt_38/if_stmt_421_if_link/if_choice_transition
      -- CP-element group 119: 	 branch_block_stmt_38/entry_bbx_xnph515
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/$entry
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_update_start_
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Sample/rr
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_38/entry_bbx_xnph515_PhiReq/$entry
      -- CP-element group 119: 	 branch_block_stmt_38/entry_bbx_xnph515_PhiReq/$exit
      -- CP-element group 119: 	 branch_block_stmt_38/merge_stmt_442_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_38/merge_stmt_442_PhiAck/$entry
      -- CP-element group 119: 	 branch_block_stmt_38/merge_stmt_442_PhiAck/$exit
      -- CP-element group 119: 	 branch_block_stmt_38/merge_stmt_442_PhiAck/dummy
      -- 
    if_choice_transition_907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_421_branch_ack_1, ack => convTranspose_CP_34_elements(119)); -- 
    rr_946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(119), ack => type_cast_457_inst_req_0); -- 
    cr_951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(119), ack => type_cast_457_inst_req_1); -- 
    -- CP-element group 120:  transition  place  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	470 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_38/if_stmt_421_else_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_38/if_stmt_421_else_link/else_choice_transition
      -- CP-element group 120: 	 branch_block_stmt_38/entry_forx_xcond190x_xpreheader
      -- CP-element group 120: 	 branch_block_stmt_38/entry_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 120: 	 branch_block_stmt_38/entry_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_421_branch_ack_0, ack => convTranspose_CP_34_elements(120)); -- 
    -- CP-element group 121:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	470 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	167 
    -- CP-element group 121: 	168 
    -- CP-element group 121:  members (18) 
      -- CP-element group 121: 	 branch_block_stmt_38/merge_stmt_643__exit__
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678__entry__
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_update_start_
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/if_stmt_436_if_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_38/if_stmt_436_if_link/if_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_38/forx_xcond190x_xpreheader_bbx_xnph511
      -- CP-element group 121: 	 branch_block_stmt_38/forx_xcond190x_xpreheader_bbx_xnph511_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/forx_xcond190x_xpreheader_bbx_xnph511_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_38/merge_stmt_643_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_38/merge_stmt_643_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/merge_stmt_643_PhiAck/$exit
      -- CP-element group 121: 	 branch_block_stmt_38/merge_stmt_643_PhiAck/dummy
      -- 
    if_choice_transition_929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_436_branch_ack_1, ack => convTranspose_CP_34_elements(121)); -- 
    cr_1310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(121), ack => type_cast_664_inst_req_1); -- 
    rr_1305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(121), ack => type_cast_664_inst_req_0); -- 
    -- CP-element group 122:  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	470 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	483 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_38/if_stmt_436_else_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_38/if_stmt_436_else_link/else_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_38/forx_xcond190x_xpreheader_forx_xend250
      -- CP-element group 122: 	 branch_block_stmt_38/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_38/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$exit
      -- 
    else_choice_transition_933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_436_branch_ack_0, ack => convTranspose_CP_34_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	119 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Sample/ra
      -- 
    ra_947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_457_inst_ack_0, ack => convTranspose_CP_34_elements(123)); -- 
    -- CP-element group 124:  transition  place  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	119 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	471 
    -- CP-element group 124:  members (9) 
      -- CP-element group 124: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471__exit__
      -- CP-element group 124: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody
      -- CP-element group 124: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/$exit
      -- CP-element group 124: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Update/ca
      -- CP-element group 124: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/$entry
      -- CP-element group 124: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_474/$entry
      -- CP-element group 124: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/$entry
      -- 
    ca_952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_457_inst_ack_1, ack => convTranspose_CP_34_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	476 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	164 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_sample_complete
      -- CP-element group 125: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Sample/ack
      -- 
    ack_981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_486_index_offset_ack_0, ack => convTranspose_CP_34_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	476 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (11) 
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_root_address_calculated
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_offset_calculated
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Update/ack
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_base_plus_offset/$entry
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_base_plus_offset/$exit
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_base_plus_offset/sum_rename_req
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_base_plus_offset/sum_rename_ack
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_request/$entry
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_request/req
      -- 
    ack_986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_486_index_offset_ack_1, ack => convTranspose_CP_34_elements(126)); -- 
    req_995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(126), ack => addr_of_487_final_reg_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_request/$exit
      -- CP-element group 127: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_request/ack
      -- 
    ack_996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_487_final_reg_ack_0, ack => convTranspose_CP_34_elements(127)); -- 
    -- CP-element group 128:  fork  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	476 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	161 
    -- CP-element group 128:  members (19) 
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_word_addrgen/root_register_ack
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_word_addrgen/root_register_req
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_word_addrgen/$exit
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_word_addrgen/$entry
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_plus_offset/sum_rename_ack
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_plus_offset/sum_rename_req
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_plus_offset/$exit
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_plus_offset/$entry
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_addr_resize/base_resize_ack
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_addr_resize/base_resize_req
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_addr_resize/$exit
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_addr_resize/$entry
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_address_resized
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_root_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_word_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_complete/$exit
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_complete/ack
      -- 
    ack_1001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_487_final_reg_ack_1, ack => convTranspose_CP_34_elements(128)); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	476 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_update_start_
      -- CP-element group 129: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Sample/ra
      -- CP-element group 129: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Update/cr
      -- 
    ra_1010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_490_inst_ack_0, ack => convTranspose_CP_34_elements(129)); -- 
    cr_1014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(129), ack => RPIPE_ConvTranspose_input_pipe_490_inst_req_1); -- 
    -- CP-element group 130:  fork  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (9) 
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Sample/rr
      -- 
    ca_1015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_490_inst_ack_1, ack => convTranspose_CP_34_elements(130)); -- 
    rr_1023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(130), ack => type_cast_494_inst_req_0); -- 
    rr_1037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(130), ack => RPIPE_ConvTranspose_input_pipe_503_inst_req_0); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Sample/ra
      -- 
    ra_1024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_494_inst_ack_0, ack => convTranspose_CP_34_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	476 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	161 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Update/ca
      -- 
    ca_1029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_494_inst_ack_1, ack => convTranspose_CP_34_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_update_start_
      -- CP-element group 133: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Update/cr
      -- 
    ra_1038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_503_inst_ack_0, ack => convTranspose_CP_34_elements(133)); -- 
    cr_1042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(133), ack => RPIPE_ConvTranspose_input_pipe_503_inst_req_1); -- 
    -- CP-element group 134:  fork  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (9) 
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Sample/rr
      -- 
    ca_1043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_503_inst_ack_1, ack => convTranspose_CP_34_elements(134)); -- 
    rr_1051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(134), ack => type_cast_507_inst_req_0); -- 
    rr_1065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(134), ack => RPIPE_ConvTranspose_input_pipe_521_inst_req_0); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Sample/ra
      -- 
    ra_1052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_507_inst_ack_0, ack => convTranspose_CP_34_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	476 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	161 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Update/ca
      -- 
    ca_1057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_507_inst_ack_1, ack => convTranspose_CP_34_elements(136)); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_update_start_
      -- CP-element group 137: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Sample/ra
      -- CP-element group 137: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Update/cr
      -- 
    ra_1066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_521_inst_ack_0, ack => convTranspose_CP_34_elements(137)); -- 
    cr_1070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(137), ack => RPIPE_ConvTranspose_input_pipe_521_inst_req_1); -- 
    -- CP-element group 138:  fork  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138: 	141 
    -- CP-element group 138:  members (9) 
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Update/ca
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Sample/rr
      -- 
    ca_1071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_521_inst_ack_1, ack => convTranspose_CP_34_elements(138)); -- 
    rr_1079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(138), ack => type_cast_525_inst_req_0); -- 
    rr_1093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(138), ack => RPIPE_ConvTranspose_input_pipe_539_inst_req_0); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Sample/ra
      -- 
    ra_1080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_525_inst_ack_0, ack => convTranspose_CP_34_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	476 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	161 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Update/ca
      -- 
    ca_1085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_525_inst_ack_1, ack => convTranspose_CP_34_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	138 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (6) 
      -- CP-element group 141: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Update/cr
      -- CP-element group 141: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Sample/ra
      -- CP-element group 141: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_update_start_
      -- CP-element group 141: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_sample_completed_
      -- 
    ra_1094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_539_inst_ack_0, ack => convTranspose_CP_34_elements(141)); -- 
    cr_1098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(141), ack => RPIPE_ConvTranspose_input_pipe_539_inst_req_1); -- 
    -- CP-element group 142:  fork  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	145 
    -- CP-element group 142:  members (9) 
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Update/ca
      -- 
    ca_1099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_539_inst_ack_1, ack => convTranspose_CP_34_elements(142)); -- 
    rr_1107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(142), ack => type_cast_543_inst_req_0); -- 
    rr_1121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(142), ack => RPIPE_ConvTranspose_input_pipe_557_inst_req_0); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_sample_completed_
      -- 
    ra_1108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_543_inst_ack_0, ack => convTranspose_CP_34_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	476 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	161 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_update_completed_
      -- 
    ca_1113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_543_inst_ack_1, ack => convTranspose_CP_34_elements(144)); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	142 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_update_start_
      -- CP-element group 145: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Sample/$exit
      -- 
    ra_1122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_557_inst_ack_0, ack => convTranspose_CP_34_elements(145)); -- 
    cr_1126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(145), ack => RPIPE_ConvTranspose_input_pipe_557_inst_req_1); -- 
    -- CP-element group 146:  fork  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	149 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Update/$exit
      -- 
    ca_1127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_557_inst_ack_1, ack => convTranspose_CP_34_elements(146)); -- 
    rr_1135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(146), ack => type_cast_561_inst_req_0); -- 
    rr_1149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(146), ack => RPIPE_ConvTranspose_input_pipe_575_inst_req_0); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_sample_completed_
      -- 
    ra_1136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_561_inst_ack_0, ack => convTranspose_CP_34_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	476 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	161 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_update_completed_
      -- 
    ca_1141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_561_inst_ack_1, ack => convTranspose_CP_34_elements(148)); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	146 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_update_start_
      -- CP-element group 149: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_sample_completed_
      -- 
    ra_1150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_575_inst_ack_0, ack => convTranspose_CP_34_elements(149)); -- 
    cr_1154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(149), ack => RPIPE_ConvTranspose_input_pipe_575_inst_req_1); -- 
    -- CP-element group 150:  fork  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (9) 
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_update_completed_
      -- 
    ca_1155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_575_inst_ack_1, ack => convTranspose_CP_34_elements(150)); -- 
    rr_1163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(150), ack => type_cast_579_inst_req_0); -- 
    rr_1177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(150), ack => RPIPE_ConvTranspose_input_pipe_593_inst_req_0); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_sample_completed_
      -- 
    ra_1164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_579_inst_ack_0, ack => convTranspose_CP_34_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	476 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	161 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_update_completed_
      -- 
    ca_1169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_579_inst_ack_1, ack => convTranspose_CP_34_elements(152)); -- 
    -- CP-element group 153:  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	150 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (6) 
      -- CP-element group 153: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Update/cr
      -- CP-element group 153: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_update_start_
      -- CP-element group 153: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_sample_completed_
      -- 
    ra_1178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_593_inst_ack_0, ack => convTranspose_CP_34_elements(153)); -- 
    cr_1182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(153), ack => RPIPE_ConvTranspose_input_pipe_593_inst_req_1); -- 
    -- CP-element group 154:  fork  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154: 	157 
    -- CP-element group 154:  members (9) 
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_sample_start_
      -- 
    ca_1183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_593_inst_ack_1, ack => convTranspose_CP_34_elements(154)); -- 
    rr_1191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(154), ack => type_cast_597_inst_req_0); -- 
    rr_1205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(154), ack => RPIPE_ConvTranspose_input_pipe_611_inst_req_0); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Sample/ra
      -- CP-element group 155: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Sample/$exit
      -- 
    ra_1192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_597_inst_ack_0, ack => convTranspose_CP_34_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	476 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	161 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Update/ca
      -- CP-element group 156: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Update/$exit
      -- 
    ca_1197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_597_inst_ack_1, ack => convTranspose_CP_34_elements(156)); -- 
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Update/cr
      -- CP-element group 157: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Sample/ra
      -- CP-element group 157: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_update_start_
      -- CP-element group 157: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_sample_completed_
      -- 
    ra_1206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_611_inst_ack_0, ack => convTranspose_CP_34_elements(157)); -- 
    cr_1210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(157), ack => RPIPE_ConvTranspose_input_pipe_611_inst_req_1); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Sample/rr
      -- CP-element group 158: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Update/ca
      -- CP-element group 158: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_update_completed_
      -- 
    ca_1211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_611_inst_ack_1, ack => convTranspose_CP_34_elements(158)); -- 
    rr_1219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(158), ack => type_cast_615_inst_req_0); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Sample/ra
      -- CP-element group 159: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_sample_completed_
      -- 
    ra_1220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_615_inst_ack_0, ack => convTranspose_CP_34_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	476 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Update/ca
      -- CP-element group 160: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_update_completed_
      -- 
    ca_1225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_615_inst_ack_1, ack => convTranspose_CP_34_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	128 
    -- CP-element group 161: 	132 
    -- CP-element group 161: 	136 
    -- CP-element group 161: 	140 
    -- CP-element group 161: 	144 
    -- CP-element group 161: 	148 
    -- CP-element group 161: 	152 
    -- CP-element group 161: 	156 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (9) 
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/word_access_start/word_0/rr
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/word_access_start/word_0/$entry
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/word_access_start/$entry
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/ptr_deref_623_Split/split_ack
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/ptr_deref_623_Split/split_req
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/ptr_deref_623_Split/$exit
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/ptr_deref_623_Split/$entry
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_sample_start_
      -- 
    rr_1263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(161), ack => ptr_deref_623_store_0_req_0); -- 
    convTranspose_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(128) & convTranspose_CP_34_elements(132) & convTranspose_CP_34_elements(136) & convTranspose_CP_34_elements(140) & convTranspose_CP_34_elements(144) & convTranspose_CP_34_elements(148) & convTranspose_CP_34_elements(152) & convTranspose_CP_34_elements(156) & convTranspose_CP_34_elements(160);
      gj_convTranspose_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/word_access_start/word_0/ra
      -- CP-element group 162: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/word_access_start/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/word_access_start/$exit
      -- CP-element group 162: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_sample_completed_
      -- 
    ra_1264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_623_store_0_ack_0, ack => convTranspose_CP_34_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	476 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/word_access_complete/$exit
      -- CP-element group 163: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/word_access_complete/word_0/ca
      -- CP-element group 163: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/word_access_complete/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_update_completed_
      -- 
    ca_1275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_623_store_0_ack_1, ack => convTranspose_CP_34_elements(163)); -- 
    -- CP-element group 164:  branch  join  transition  place  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: 	125 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (10) 
      -- CP-element group 164: 	 branch_block_stmt_38/if_stmt_637_eval_test/$exit
      -- CP-element group 164: 	 branch_block_stmt_38/if_stmt_637_eval_test/branch_req
      -- CP-element group 164: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636__exit__
      -- CP-element group 164: 	 branch_block_stmt_38/if_stmt_637__entry__
      -- CP-element group 164: 	 branch_block_stmt_38/if_stmt_637_eval_test/$entry
      -- CP-element group 164: 	 branch_block_stmt_38/if_stmt_637_dead_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_38/R_exitcond3_638_place
      -- CP-element group 164: 	 branch_block_stmt_38/if_stmt_637_else_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_38/if_stmt_637_if_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/$exit
      -- 
    branch_req_1283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(164), ack => if_stmt_637_branch_req_0); -- 
    convTranspose_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(163) & convTranspose_CP_34_elements(125);
      gj_convTranspose_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  merge  transition  place  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	470 
    -- CP-element group 165:  members (13) 
      -- CP-element group 165: 	 branch_block_stmt_38/merge_stmt_427__exit__
      -- CP-element group 165: 	 branch_block_stmt_38/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader
      -- CP-element group 165: 	 branch_block_stmt_38/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit
      -- CP-element group 165: 	 branch_block_stmt_38/if_stmt_637_if_link/if_choice_transition
      -- CP-element group 165: 	 branch_block_stmt_38/if_stmt_637_if_link/$exit
      -- CP-element group 165: 	 branch_block_stmt_38/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_38/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_38/merge_stmt_427_PhiReqMerge
      -- CP-element group 165: 	 branch_block_stmt_38/merge_stmt_427_PhiAck/$entry
      -- CP-element group 165: 	 branch_block_stmt_38/merge_stmt_427_PhiAck/$exit
      -- CP-element group 165: 	 branch_block_stmt_38/merge_stmt_427_PhiAck/dummy
      -- CP-element group 165: 	 branch_block_stmt_38/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_38/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_637_branch_ack_1, ack => convTranspose_CP_34_elements(165)); -- 
    -- CP-element group 166:  fork  transition  place  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	472 
    -- CP-element group 166: 	473 
    -- CP-element group 166:  members (12) 
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody
      -- CP-element group 166: 	 branch_block_stmt_38/if_stmt_637_else_link/else_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_38/if_stmt_637_else_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/$entry
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/$entry
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/$entry
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/$entry
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_637_branch_ack_0, ack => convTranspose_CP_34_elements(166)); -- 
    rr_3511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(166), ack => type_cast_480_inst_req_0); -- 
    cr_3516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(166), ack => type_cast_480_inst_req_1); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	121 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Sample/ra
      -- CP-element group 167: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_sample_completed_
      -- 
    ra_1306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_664_inst_ack_0, ack => convTranspose_CP_34_elements(167)); -- 
    -- CP-element group 168:  transition  place  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	121 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	477 
    -- CP-element group 168:  members (9) 
      -- CP-element group 168: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678__exit__
      -- CP-element group 168: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196
      -- CP-element group 168: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Update/ca
      -- CP-element group 168: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/$exit
      -- CP-element group 168: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/$entry
      -- CP-element group 168: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_681/$entry
      -- CP-element group 168: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/$entry
      -- 
    ca_1311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_664_inst_ack_1, ack => convTranspose_CP_34_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	482 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	208 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Sample/ack
      -- CP-element group 169: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_sample_complete
      -- 
    ack_1340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_693_index_offset_ack_0, ack => convTranspose_CP_34_elements(169)); -- 
    -- CP-element group 170:  transition  input  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	482 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (11) 
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_request/req
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_request/$entry
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_base_plus_offset/$entry
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_base_plus_offset/sum_rename_ack
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_base_plus_offset/sum_rename_req
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_base_plus_offset/$exit
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_offset_calculated
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_root_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Update/ack
      -- 
    ack_1345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_693_index_offset_ack_1, ack => convTranspose_CP_34_elements(170)); -- 
    req_1354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(170), ack => addr_of_694_final_reg_req_0); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_request/$exit
      -- CP-element group 171: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_request/ack
      -- 
    ack_1355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_694_final_reg_ack_0, ack => convTranspose_CP_34_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	482 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	205 
    -- CP-element group 172:  members (19) 
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_complete/ack
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_complete/$exit
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_word_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_address_resized
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_addr_resize/$entry
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_addr_resize/$exit
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_addr_resize/base_resize_req
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_addr_resize/base_resize_ack
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_word_addrgen/$entry
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_word_addrgen/$exit
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_word_addrgen/root_register_req
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_word_addrgen/root_register_ack
      -- 
    ack_1360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_694_final_reg_ack_1, ack => convTranspose_CP_34_elements(172)); -- 
    -- CP-element group 173:  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	482 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Update/cr
      -- CP-element group 173: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Sample/ra
      -- CP-element group 173: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_update_start_
      -- CP-element group 173: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_sample_completed_
      -- 
    ra_1369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_697_inst_ack_0, ack => convTranspose_CP_34_elements(173)); -- 
    cr_1373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(173), ack => RPIPE_ConvTranspose_input_pipe_697_inst_req_1); -- 
    -- CP-element group 174:  fork  transition  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174: 	177 
    -- CP-element group 174:  members (9) 
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Update/ca
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Sample/$entry
      -- 
    ca_1374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_697_inst_ack_1, ack => convTranspose_CP_34_elements(174)); -- 
    rr_1382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(174), ack => type_cast_701_inst_req_0); -- 
    rr_1396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(174), ack => RPIPE_ConvTranspose_input_pipe_710_inst_req_0); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Sample/$exit
      -- 
    ra_1383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_701_inst_ack_0, ack => convTranspose_CP_34_elements(175)); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	482 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	205 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_update_completed_
      -- 
    ca_1388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_701_inst_ack_1, ack => convTranspose_CP_34_elements(176)); -- 
    -- CP-element group 177:  transition  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	174 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (6) 
      -- CP-element group 177: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_update_start_
      -- 
    ra_1397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_710_inst_ack_0, ack => convTranspose_CP_34_elements(177)); -- 
    cr_1401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(177), ack => RPIPE_ConvTranspose_input_pipe_710_inst_req_1); -- 
    -- CP-element group 178:  fork  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178: 	181 
    -- CP-element group 178:  members (9) 
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Sample/$entry
      -- 
    ca_1402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_710_inst_ack_1, ack => convTranspose_CP_34_elements(178)); -- 
    rr_1410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(178), ack => type_cast_714_inst_req_0); -- 
    rr_1424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(178), ack => RPIPE_ConvTranspose_input_pipe_728_inst_req_0); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_sample_completed_
      -- 
    ra_1411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_714_inst_ack_0, ack => convTranspose_CP_34_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	482 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	205 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_update_completed_
      -- 
    ca_1416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_714_inst_ack_1, ack => convTranspose_CP_34_elements(180)); -- 
    -- CP-element group 181:  transition  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	178 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (6) 
      -- CP-element group 181: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_update_start_
      -- CP-element group 181: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Update/cr
      -- CP-element group 181: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Sample/ra
      -- CP-element group 181: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Sample/$exit
      -- 
    ra_1425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_728_inst_ack_0, ack => convTranspose_CP_34_elements(181)); -- 
    cr_1429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(181), ack => RPIPE_ConvTranspose_input_pipe_728_inst_req_1); -- 
    -- CP-element group 182:  fork  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182: 	185 
    -- CP-element group 182:  members (9) 
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Update/ca
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_update_completed_
      -- 
    ca_1430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_728_inst_ack_1, ack => convTranspose_CP_34_elements(182)); -- 
    rr_1438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(182), ack => type_cast_732_inst_req_0); -- 
    rr_1452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(182), ack => RPIPE_ConvTranspose_input_pipe_746_inst_req_0); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Sample/ra
      -- 
    ra_1439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_732_inst_ack_0, ack => convTranspose_CP_34_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	482 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	205 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Update/$exit
      -- 
    ca_1444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_732_inst_ack_1, ack => convTranspose_CP_34_elements(184)); -- 
    -- CP-element group 185:  transition  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	182 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (6) 
      -- CP-element group 185: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Update/cr
      -- CP-element group 185: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Sample/ra
      -- CP-element group 185: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_update_start_
      -- CP-element group 185: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_sample_completed_
      -- 
    ra_1453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_746_inst_ack_0, ack => convTranspose_CP_34_elements(185)); -- 
    cr_1457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(185), ack => RPIPE_ConvTranspose_input_pipe_746_inst_req_1); -- 
    -- CP-element group 186:  fork  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	189 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (9) 
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Update/ca
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Sample/rr
      -- 
    ca_1458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_746_inst_ack_1, ack => convTranspose_CP_34_elements(186)); -- 
    rr_1480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(186), ack => RPIPE_ConvTranspose_input_pipe_764_inst_req_0); -- 
    rr_1466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(186), ack => type_cast_750_inst_req_0); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Sample/ra
      -- 
    ra_1467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_750_inst_ack_0, ack => convTranspose_CP_34_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	482 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	205 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Update/ca
      -- 
    ca_1472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_750_inst_ack_1, ack => convTranspose_CP_34_elements(188)); -- 
    -- CP-element group 189:  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	186 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (6) 
      -- CP-element group 189: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_update_start_
      -- CP-element group 189: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Update/cr
      -- 
    ra_1481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_764_inst_ack_0, ack => convTranspose_CP_34_elements(189)); -- 
    cr_1485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(189), ack => RPIPE_ConvTranspose_input_pipe_764_inst_req_1); -- 
    -- CP-element group 190:  fork  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	193 
    -- CP-element group 190: 	191 
    -- CP-element group 190:  members (9) 
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Sample/rr
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Sample/rr
      -- 
    ca_1486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_764_inst_ack_1, ack => convTranspose_CP_34_elements(190)); -- 
    rr_1494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(190), ack => type_cast_768_inst_req_0); -- 
    rr_1508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(190), ack => RPIPE_ConvTranspose_input_pipe_782_inst_req_0); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Sample/ra
      -- 
    ra_1495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_768_inst_ack_0, ack => convTranspose_CP_34_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	482 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	205 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Update/ca
      -- 
    ca_1500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_768_inst_ack_1, ack => convTranspose_CP_34_elements(192)); -- 
    -- CP-element group 193:  transition  input  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	190 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (6) 
      -- CP-element group 193: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_update_start_
      -- CP-element group 193: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Sample/ra
      -- CP-element group 193: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Update/$entry
      -- CP-element group 193: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Update/cr
      -- 
    ra_1509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_782_inst_ack_0, ack => convTranspose_CP_34_elements(193)); -- 
    cr_1513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(193), ack => RPIPE_ConvTranspose_input_pipe_782_inst_req_1); -- 
    -- CP-element group 194:  fork  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: 	197 
    -- CP-element group 194:  members (9) 
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Sample/rr
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Sample/rr
      -- 
    ca_1514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_782_inst_ack_1, ack => convTranspose_CP_34_elements(194)); -- 
    rr_1522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(194), ack => type_cast_786_inst_req_0); -- 
    rr_1536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(194), ack => RPIPE_ConvTranspose_input_pipe_800_inst_req_0); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Sample/ra
      -- 
    ra_1523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_786_inst_ack_0, ack => convTranspose_CP_34_elements(195)); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	482 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	205 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Update/ca
      -- 
    ca_1528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_786_inst_ack_1, ack => convTranspose_CP_34_elements(196)); -- 
    -- CP-element group 197:  transition  input  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	194 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (6) 
      -- CP-element group 197: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_update_start_
      -- CP-element group 197: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Sample/ra
      -- CP-element group 197: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Update/cr
      -- 
    ra_1537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_800_inst_ack_0, ack => convTranspose_CP_34_elements(197)); -- 
    cr_1541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(197), ack => RPIPE_ConvTranspose_input_pipe_800_inst_req_1); -- 
    -- CP-element group 198:  fork  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198: 	201 
    -- CP-element group 198:  members (9) 
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Update/ca
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Sample/rr
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Sample/rr
      -- 
    ca_1542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_800_inst_ack_1, ack => convTranspose_CP_34_elements(198)); -- 
    rr_1550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(198), ack => type_cast_804_inst_req_0); -- 
    rr_1564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(198), ack => RPIPE_ConvTranspose_input_pipe_818_inst_req_0); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Sample/ra
      -- 
    ra_1551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_804_inst_ack_0, ack => convTranspose_CP_34_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	482 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	205 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Update/ca
      -- 
    ca_1556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_804_inst_ack_1, ack => convTranspose_CP_34_elements(200)); -- 
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	198 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_update_start_
      -- CP-element group 201: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Sample/ra
      -- CP-element group 201: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Update/cr
      -- 
    ra_1565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_818_inst_ack_0, ack => convTranspose_CP_34_elements(201)); -- 
    cr_1569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(201), ack => RPIPE_ConvTranspose_input_pipe_818_inst_req_1); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Update/ca
      -- CP-element group 202: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Sample/rr
      -- 
    ca_1570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_818_inst_ack_1, ack => convTranspose_CP_34_elements(202)); -- 
    rr_1578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(202), ack => type_cast_822_inst_req_0); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Sample/ra
      -- 
    ra_1579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_822_inst_ack_0, ack => convTranspose_CP_34_elements(203)); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	482 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Update/ca
      -- 
    ca_1584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_822_inst_ack_1, ack => convTranspose_CP_34_elements(204)); -- 
    -- CP-element group 205:  join  transition  output  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	196 
    -- CP-element group 205: 	200 
    -- CP-element group 205: 	204 
    -- CP-element group 205: 	188 
    -- CP-element group 205: 	192 
    -- CP-element group 205: 	172 
    -- CP-element group 205: 	176 
    -- CP-element group 205: 	180 
    -- CP-element group 205: 	184 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (9) 
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_sample_start_
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/$entry
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/ptr_deref_830_Split/$entry
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/ptr_deref_830_Split/$exit
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/ptr_deref_830_Split/split_req
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/ptr_deref_830_Split/split_ack
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/word_access_start/$entry
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/word_access_start/word_0/$entry
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/word_access_start/word_0/rr
      -- 
    rr_1622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(205), ack => ptr_deref_830_store_0_req_0); -- 
    convTranspose_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(196) & convTranspose_CP_34_elements(200) & convTranspose_CP_34_elements(204) & convTranspose_CP_34_elements(188) & convTranspose_CP_34_elements(192) & convTranspose_CP_34_elements(172) & convTranspose_CP_34_elements(176) & convTranspose_CP_34_elements(180) & convTranspose_CP_34_elements(184);
      gj_convTranspose_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (5) 
      -- CP-element group 206: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_sample_completed_
      -- CP-element group 206: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/word_access_start/$exit
      -- CP-element group 206: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/word_access_start/word_0/$exit
      -- CP-element group 206: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/word_access_start/word_0/ra
      -- 
    ra_1623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_830_store_0_ack_0, ack => convTranspose_CP_34_elements(206)); -- 
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	482 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (5) 
      -- CP-element group 207: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_update_completed_
      -- CP-element group 207: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/word_access_complete/$exit
      -- CP-element group 207: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/word_access_complete/word_0/$exit
      -- CP-element group 207: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/word_access_complete/word_0/ca
      -- 
    ca_1634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_830_store_0_ack_1, ack => convTranspose_CP_34_elements(207)); -- 
    -- CP-element group 208:  branch  join  transition  place  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: 	169 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (10) 
      -- CP-element group 208: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843__exit__
      -- CP-element group 208: 	 branch_block_stmt_38/if_stmt_844__entry__
      -- CP-element group 208: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/$exit
      -- CP-element group 208: 	 branch_block_stmt_38/if_stmt_844_dead_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_38/if_stmt_844_eval_test/$entry
      -- CP-element group 208: 	 branch_block_stmt_38/if_stmt_844_eval_test/$exit
      -- CP-element group 208: 	 branch_block_stmt_38/if_stmt_844_eval_test/branch_req
      -- CP-element group 208: 	 branch_block_stmt_38/R_exitcond2_845_place
      -- CP-element group 208: 	 branch_block_stmt_38/if_stmt_844_if_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_38/if_stmt_844_else_link/$entry
      -- 
    branch_req_1642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(208), ack => if_stmt_844_branch_req_0); -- 
    convTranspose_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(207) & convTranspose_CP_34_elements(169);
      gj_convTranspose_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  merge  transition  place  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	483 
    -- CP-element group 209:  members (13) 
      -- CP-element group 209: 	 branch_block_stmt_38/merge_stmt_850__exit__
      -- CP-element group 209: 	 branch_block_stmt_38/forx_xend250x_xloopexit_forx_xend250
      -- CP-element group 209: 	 branch_block_stmt_38/if_stmt_844_if_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_38/if_stmt_844_if_link/if_choice_transition
      -- CP-element group 209: 	 branch_block_stmt_38/forx_xbody196_forx_xend250x_xloopexit
      -- CP-element group 209: 	 branch_block_stmt_38/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_38/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$exit
      -- CP-element group 209: 	 branch_block_stmt_38/merge_stmt_850_PhiReqMerge
      -- CP-element group 209: 	 branch_block_stmt_38/merge_stmt_850_PhiAck/$entry
      -- CP-element group 209: 	 branch_block_stmt_38/merge_stmt_850_PhiAck/$exit
      -- CP-element group 209: 	 branch_block_stmt_38/merge_stmt_850_PhiAck/dummy
      -- CP-element group 209: 	 branch_block_stmt_38/forx_xend250x_xloopexit_forx_xend250_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_38/forx_xend250x_xloopexit_forx_xend250_PhiReq/$exit
      -- 
    if_choice_transition_1647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_844_branch_ack_1, ack => convTranspose_CP_34_elements(209)); -- 
    -- CP-element group 210:  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	478 
    -- CP-element group 210: 	479 
    -- CP-element group 210:  members (12) 
      -- CP-element group 210: 	 branch_block_stmt_38/if_stmt_844_else_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_38/if_stmt_844_else_link/else_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/$entry
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/$entry
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_844_branch_ack_0, ack => convTranspose_CP_34_elements(210)); -- 
    rr_3565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(210), ack => type_cast_687_inst_req_0); -- 
    cr_3570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(210), ack => type_cast_687_inst_req_1); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	483 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Sample/ra
      -- 
    ra_1665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_855_inst_ack_0, ack => convTranspose_CP_34_elements(211)); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	483 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	217 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Update/ca
      -- 
    ca_1670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_855_inst_ack_1, ack => convTranspose_CP_34_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	483 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Sample/ra
      -- 
    ra_1679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_859_inst_ack_0, ack => convTranspose_CP_34_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	483 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	217 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Update/ca
      -- 
    ca_1684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_859_inst_ack_1, ack => convTranspose_CP_34_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	483 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Sample/ra
      -- 
    ra_1693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_863_inst_ack_0, ack => convTranspose_CP_34_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	483 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Update/ca
      -- 
    ca_1698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_863_inst_ack_1, ack => convTranspose_CP_34_elements(216)); -- 
    -- CP-element group 217:  branch  join  transition  place  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	212 
    -- CP-element group 217: 	214 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (10) 
      -- CP-element group 217: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880__exit__
      -- CP-element group 217: 	 branch_block_stmt_38/if_stmt_881__entry__
      -- CP-element group 217: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/$exit
      -- CP-element group 217: 	 branch_block_stmt_38/if_stmt_881_dead_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_38/if_stmt_881_eval_test/$entry
      -- CP-element group 217: 	 branch_block_stmt_38/if_stmt_881_eval_test/$exit
      -- CP-element group 217: 	 branch_block_stmt_38/if_stmt_881_eval_test/branch_req
      -- CP-element group 217: 	 branch_block_stmt_38/R_cmp264505_882_place
      -- CP-element group 217: 	 branch_block_stmt_38/if_stmt_881_if_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_38/if_stmt_881_else_link/$entry
      -- 
    branch_req_1706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(217), ack => if_stmt_881_branch_req_0); -- 
    convTranspose_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(212) & convTranspose_CP_34_elements(214) & convTranspose_CP_34_elements(216);
      gj_convTranspose_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: 	221 
    -- CP-element group 218:  members (18) 
      -- CP-element group 218: 	 branch_block_stmt_38/merge_stmt_887__exit__
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922__entry__
      -- CP-element group 218: 	 branch_block_stmt_38/if_stmt_881_if_link/$exit
      -- CP-element group 218: 	 branch_block_stmt_38/if_stmt_881_if_link/if_choice_transition
      -- CP-element group 218: 	 branch_block_stmt_38/forx_xend250_bbx_xnph507
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/$entry
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_update_start_
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Sample/rr
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_38/forx_xend250_bbx_xnph507_PhiReq/$entry
      -- CP-element group 218: 	 branch_block_stmt_38/forx_xend250_bbx_xnph507_PhiReq/$exit
      -- CP-element group 218: 	 branch_block_stmt_38/merge_stmt_887_PhiReqMerge
      -- CP-element group 218: 	 branch_block_stmt_38/merge_stmt_887_PhiAck/$entry
      -- CP-element group 218: 	 branch_block_stmt_38/merge_stmt_887_PhiAck/$exit
      -- CP-element group 218: 	 branch_block_stmt_38/merge_stmt_887_PhiAck/dummy
      -- 
    if_choice_transition_1711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_881_branch_ack_1, ack => convTranspose_CP_34_elements(218)); -- 
    rr_1728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(218), ack => type_cast_908_inst_req_0); -- 
    cr_1733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(218), ack => type_cast_908_inst_req_1); -- 
    -- CP-element group 219:  transition  place  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	490 
    -- CP-element group 219:  members (5) 
      -- CP-element group 219: 	 branch_block_stmt_38/if_stmt_881_else_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_38/if_stmt_881_else_link/else_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_38/forx_xend250_forx_xend273
      -- CP-element group 219: 	 branch_block_stmt_38/forx_xend250_forx_xend273_PhiReq/$entry
      -- CP-element group 219: 	 branch_block_stmt_38/forx_xend250_forx_xend273_PhiReq/$exit
      -- 
    else_choice_transition_1715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_881_branch_ack_0, ack => convTranspose_CP_34_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Sample/ra
      -- 
    ra_1729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_908_inst_ack_0, ack => convTranspose_CP_34_elements(220)); -- 
    -- CP-element group 221:  transition  place  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	218 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	484 
    -- CP-element group 221:  members (9) 
      -- CP-element group 221: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922__exit__
      -- CP-element group 221: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266
      -- CP-element group 221: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/$exit
      -- CP-element group 221: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Update/ca
      -- CP-element group 221: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_925/$entry
      -- CP-element group 221: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/$entry
      -- 
    ca_1734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_908_inst_ack_1, ack => convTranspose_CP_34_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	489 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	228 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_sample_complete
      -- CP-element group 222: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Sample/ack
      -- 
    ack_1763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_937_index_offset_ack_0, ack => convTranspose_CP_34_elements(222)); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	489 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (11) 
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_root_address_calculated
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_offset_calculated
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Update/ack
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_base_plus_offset/$entry
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_base_plus_offset/$exit
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_base_plus_offset/sum_rename_req
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_base_plus_offset/sum_rename_ack
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_request/$entry
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_request/req
      -- 
    ack_1768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_937_index_offset_ack_1, ack => convTranspose_CP_34_elements(223)); -- 
    req_1777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(223), ack => addr_of_938_final_reg_req_0); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_request/$exit
      -- CP-element group 224: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_request/ack
      -- 
    ack_1778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_938_final_reg_ack_0, ack => convTranspose_CP_34_elements(224)); -- 
    -- CP-element group 225:  join  fork  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	489 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (28) 
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_complete/$exit
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_complete/ack
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_word_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_root_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_address_resized
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_addr_resize/$entry
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_addr_resize/$exit
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_addr_resize/base_resize_req
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_addr_resize/base_resize_ack
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_plus_offset/$entry
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_plus_offset/$exit
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_plus_offset/sum_rename_req
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_plus_offset/sum_rename_ack
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_word_addrgen/$entry
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_word_addrgen/$exit
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_word_addrgen/root_register_req
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_word_addrgen/root_register_ack
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/ptr_deref_941_Split/$entry
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/ptr_deref_941_Split/$exit
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/ptr_deref_941_Split/split_req
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/ptr_deref_941_Split/split_ack
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/word_access_start/$entry
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/word_access_start/word_0/$entry
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/word_access_start/word_0/rr
      -- 
    ack_1783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_938_final_reg_ack_1, ack => convTranspose_CP_34_elements(225)); -- 
    rr_1821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(225), ack => ptr_deref_941_store_0_req_0); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (5) 
      -- CP-element group 226: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/word_access_start/$exit
      -- CP-element group 226: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/word_access_start/word_0/$exit
      -- CP-element group 226: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/word_access_start/word_0/ra
      -- 
    ra_1822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_941_store_0_ack_0, ack => convTranspose_CP_34_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	489 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/word_access_complete/$exit
      -- CP-element group 227: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/word_access_complete/word_0/$exit
      -- CP-element group 227: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/word_access_complete/word_0/ca
      -- 
    ca_1833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_941_store_0_ack_1, ack => convTranspose_CP_34_elements(227)); -- 
    -- CP-element group 228:  branch  join  transition  place  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	227 
    -- CP-element group 228: 	222 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (10) 
      -- CP-element group 228: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955__exit__
      -- CP-element group 228: 	 branch_block_stmt_38/if_stmt_956__entry__
      -- CP-element group 228: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/$exit
      -- CP-element group 228: 	 branch_block_stmt_38/if_stmt_956_dead_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_38/if_stmt_956_eval_test/$entry
      -- CP-element group 228: 	 branch_block_stmt_38/if_stmt_956_eval_test/$exit
      -- CP-element group 228: 	 branch_block_stmt_38/if_stmt_956_eval_test/branch_req
      -- CP-element group 228: 	 branch_block_stmt_38/R_exitcond_957_place
      -- CP-element group 228: 	 branch_block_stmt_38/if_stmt_956_if_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_38/if_stmt_956_else_link/$entry
      -- 
    branch_req_1841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(228), ack => if_stmt_956_branch_req_0); -- 
    convTranspose_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(227) & convTranspose_CP_34_elements(222);
      gj_convTranspose_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  merge  transition  place  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	490 
    -- CP-element group 229:  members (13) 
      -- CP-element group 229: 	 branch_block_stmt_38/merge_stmt_962__exit__
      -- CP-element group 229: 	 branch_block_stmt_38/forx_xend273x_xloopexit_forx_xend273
      -- CP-element group 229: 	 branch_block_stmt_38/if_stmt_956_if_link/$exit
      -- CP-element group 229: 	 branch_block_stmt_38/if_stmt_956_if_link/if_choice_transition
      -- CP-element group 229: 	 branch_block_stmt_38/forx_xbody266_forx_xend273x_xloopexit
      -- CP-element group 229: 	 branch_block_stmt_38/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_38/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$exit
      -- CP-element group 229: 	 branch_block_stmt_38/merge_stmt_962_PhiReqMerge
      -- CP-element group 229: 	 branch_block_stmt_38/merge_stmt_962_PhiAck/$entry
      -- CP-element group 229: 	 branch_block_stmt_38/merge_stmt_962_PhiAck/$exit
      -- CP-element group 229: 	 branch_block_stmt_38/merge_stmt_962_PhiAck/dummy
      -- CP-element group 229: 	 branch_block_stmt_38/forx_xend273x_xloopexit_forx_xend273_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_38/forx_xend273x_xloopexit_forx_xend273_PhiReq/$exit
      -- 
    if_choice_transition_1846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_956_branch_ack_1, ack => convTranspose_CP_34_elements(229)); -- 
    -- CP-element group 230:  fork  transition  place  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	485 
    -- CP-element group 230: 	486 
    -- CP-element group 230:  members (12) 
      -- CP-element group 230: 	 branch_block_stmt_38/if_stmt_956_else_link/$exit
      -- CP-element group 230: 	 branch_block_stmt_38/if_stmt_956_else_link/else_choice_transition
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/$entry
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/$entry
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/$entry
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/$entry
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/$entry
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Sample/rr
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_956_branch_ack_0, ack => convTranspose_CP_34_elements(230)); -- 
    rr_3642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(230), ack => type_cast_928_inst_req_0); -- 
    cr_3647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(230), ack => type_cast_928_inst_req_1); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	490 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Sample/cra
      -- 
    cra_1864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_967_call_ack_0, ack => convTranspose_CP_34_elements(231)); -- 
    -- CP-element group 232:  transition  input  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	490 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (6) 
      -- CP-element group 232: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Update/cca
      -- CP-element group 232: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Sample/rr
      -- 
    cca_1869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_967_call_ack_1, ack => convTranspose_CP_34_elements(232)); -- 
    rr_1877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(232), ack => type_cast_972_inst_req_0); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Sample/ra
      -- 
    ra_1878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_972_inst_ack_0, ack => convTranspose_CP_34_elements(233)); -- 
    -- CP-element group 234:  fork  transition  place  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	490 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	350 
    -- CP-element group 234: 	354 
    -- CP-element group 234: 	355 
    -- CP-element group 234: 	235 
    -- CP-element group 234: 	263 
    -- CP-element group 234: 	281 
    -- CP-element group 234: 	282 
    -- CP-element group 234: 	286 
    -- CP-element group 234: 	287 
    -- CP-element group 234: 	297 
    -- CP-element group 234: 	315 
    -- CP-element group 234: 	316 
    -- CP-element group 234: 	320 
    -- CP-element group 234: 	321 
    -- CP-element group 234: 	331 
    -- CP-element group 234: 	349 
    -- CP-element group 234:  members (55) 
      -- CP-element group 234: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973__exit__
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186__entry__
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_update_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_update_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/$exit
      -- CP-element group 234: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Update/ca
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_update_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_update_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_update_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_update_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_Update/cr
      -- 
    ca_1883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_972_inst_ack_1, ack => convTranspose_CP_34_elements(234)); -- 
    req_2090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => WPIPE_Block1_start_1019_inst_req_0); -- 
    cr_2221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1054_inst_req_1); -- 
    rr_2216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1054_inst_req_0); -- 
    req_2314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => WPIPE_Block2_start_1075_inst_req_0); -- 
    cr_2249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1061_inst_req_1); -- 
    rr_2244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1061_inst_req_0); -- 
    req_1894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => WPIPE_Block0_start_975_inst_req_0); -- 
    rr_2440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1110_inst_req_0); -- 
    cr_2445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1110_inst_req_1); -- 
    rr_2468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1117_inst_req_0); -- 
    cr_2473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1117_inst_req_1); -- 
    req_2538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => WPIPE_Block3_start_1131_inst_req_0); -- 
    rr_2664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1166_inst_req_0); -- 
    cr_2669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1166_inst_req_1); -- 
    rr_2692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1173_inst_req_0); -- 
    cr_2697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1173_inst_req_1); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_update_start_
      -- CP-element group 235: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_Update/req
      -- 
    ack_1895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_975_inst_ack_0, ack => convTranspose_CP_34_elements(235)); -- 
    req_1899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(235), ack => WPIPE_Block0_start_975_inst_req_1); -- 
    -- CP-element group 236:  transition  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_Sample/req
      -- CP-element group 236: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_Update/ack
      -- CP-element group 236: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_sample_start_
      -- 
    ack_1900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_975_inst_ack_1, ack => convTranspose_CP_34_elements(236)); -- 
    req_1908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(236), ack => WPIPE_Block0_start_978_inst_req_0); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_Update/req
      -- CP-element group 237: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_update_start_
      -- CP-element group 237: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_sample_completed_
      -- 
    ack_1909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_978_inst_ack_0, ack => convTranspose_CP_34_elements(237)); -- 
    req_1913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(237), ack => WPIPE_Block0_start_978_inst_req_1); -- 
    -- CP-element group 238:  transition  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_Update/ack
      -- CP-element group 238: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_Sample/req
      -- CP-element group 238: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_update_completed_
      -- 
    ack_1914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_978_inst_ack_1, ack => convTranspose_CP_34_elements(238)); -- 
    req_1922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(238), ack => WPIPE_Block0_start_981_inst_req_0); -- 
    -- CP-element group 239:  transition  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_update_start_
      -- CP-element group 239: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_Sample/ack
      -- CP-element group 239: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_Update/req
      -- 
    ack_1923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_981_inst_ack_0, ack => convTranspose_CP_34_elements(239)); -- 
    req_1927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(239), ack => WPIPE_Block0_start_981_inst_req_1); -- 
    -- CP-element group 240:  transition  input  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (6) 
      -- CP-element group 240: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_Sample/req
      -- CP-element group 240: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_sample_start_
      -- CP-element group 240: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_Update/ack
      -- CP-element group 240: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_Update/$exit
      -- 
    ack_1928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_981_inst_ack_1, ack => convTranspose_CP_34_elements(240)); -- 
    req_1936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(240), ack => WPIPE_Block0_start_984_inst_req_0); -- 
    -- CP-element group 241:  transition  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_Update/req
      -- CP-element group 241: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_Sample/ack
      -- CP-element group 241: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_update_start_
      -- CP-element group 241: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_sample_completed_
      -- 
    ack_1937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_984_inst_ack_0, ack => convTranspose_CP_34_elements(241)); -- 
    req_1941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(241), ack => WPIPE_Block0_start_984_inst_req_1); -- 
    -- CP-element group 242:  transition  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (6) 
      -- CP-element group 242: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_Update/ack
      -- CP-element group 242: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_Sample/req
      -- CP-element group 242: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_update_completed_
      -- 
    ack_1942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_984_inst_ack_1, ack => convTranspose_CP_34_elements(242)); -- 
    req_1950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(242), ack => WPIPE_Block0_start_987_inst_req_0); -- 
    -- CP-element group 243:  transition  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (6) 
      -- CP-element group 243: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_update_start_
      -- CP-element group 243: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_Update/req
      -- CP-element group 243: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_Sample/ack
      -- CP-element group 243: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_Sample/$exit
      -- 
    ack_1951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_987_inst_ack_0, ack => convTranspose_CP_34_elements(243)); -- 
    req_1955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(243), ack => WPIPE_Block0_start_987_inst_req_1); -- 
    -- CP-element group 244:  transition  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_Update/ack
      -- CP-element group 244: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_Sample/req
      -- CP-element group 244: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_Sample/$entry
      -- 
    ack_1956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_987_inst_ack_1, ack => convTranspose_CP_34_elements(244)); -- 
    req_1964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(244), ack => WPIPE_Block0_start_990_inst_req_0); -- 
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_sample_completed_
      -- CP-element group 245: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_update_start_
      -- CP-element group 245: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_Update/req
      -- CP-element group 245: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_Sample/ack
      -- CP-element group 245: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_Sample/$exit
      -- 
    ack_1965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_990_inst_ack_0, ack => convTranspose_CP_34_elements(245)); -- 
    req_1969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(245), ack => WPIPE_Block0_start_990_inst_req_1); -- 
    -- CP-element group 246:  transition  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (6) 
      -- CP-element group 246: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_Sample/req
      -- CP-element group 246: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_Update/ack
      -- CP-element group 246: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_update_completed_
      -- 
    ack_1970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_990_inst_ack_1, ack => convTranspose_CP_34_elements(246)); -- 
    req_1978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(246), ack => WPIPE_Block0_start_993_inst_req_0); -- 
    -- CP-element group 247:  transition  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_Update/req
      -- CP-element group 247: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_Sample/ack
      -- CP-element group 247: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_update_start_
      -- CP-element group 247: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_sample_completed_
      -- 
    ack_1979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_993_inst_ack_0, ack => convTranspose_CP_34_elements(247)); -- 
    req_1983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(247), ack => WPIPE_Block0_start_993_inst_req_1); -- 
    -- CP-element group 248:  transition  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (6) 
      -- CP-element group 248: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_Update/ack
      -- CP-element group 248: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_Sample/$entry
      -- CP-element group 248: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_Sample/req
      -- 
    ack_1984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_993_inst_ack_1, ack => convTranspose_CP_34_elements(248)); -- 
    req_1992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(248), ack => WPIPE_Block0_start_996_inst_req_0); -- 
    -- CP-element group 249:  transition  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (6) 
      -- CP-element group 249: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_sample_completed_
      -- CP-element group 249: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_update_start_
      -- CP-element group 249: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_Sample/ack
      -- CP-element group 249: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_Update/req
      -- 
    ack_1993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_996_inst_ack_0, ack => convTranspose_CP_34_elements(249)); -- 
    req_1997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(249), ack => WPIPE_Block0_start_996_inst_req_1); -- 
    -- CP-element group 250:  transition  input  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (6) 
      -- CP-element group 250: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_update_completed_
      -- CP-element group 250: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_Update/ack
      -- CP-element group 250: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_Sample/req
      -- 
    ack_1998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_996_inst_ack_1, ack => convTranspose_CP_34_elements(250)); -- 
    req_2006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(250), ack => WPIPE_Block0_start_999_inst_req_0); -- 
    -- CP-element group 251:  transition  input  output  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (6) 
      -- CP-element group 251: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_update_start_
      -- CP-element group 251: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_Update/req
      -- CP-element group 251: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_Sample/ack
      -- CP-element group 251: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_Sample/$exit
      -- 
    ack_2007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_999_inst_ack_0, ack => convTranspose_CP_34_elements(251)); -- 
    req_2011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(251), ack => WPIPE_Block0_start_999_inst_req_1); -- 
    -- CP-element group 252:  transition  input  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (6) 
      -- CP-element group 252: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_Sample/req
      -- CP-element group 252: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_Update/ack
      -- CP-element group 252: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_Update/$exit
      -- 
    ack_2012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_999_inst_ack_1, ack => convTranspose_CP_34_elements(252)); -- 
    req_2020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(252), ack => WPIPE_Block0_start_1002_inst_req_0); -- 
    -- CP-element group 253:  transition  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (6) 
      -- CP-element group 253: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_Sample/ack
      -- CP-element group 253: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_update_start_
      -- CP-element group 253: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_Update/req
      -- CP-element group 253: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_sample_completed_
      -- 
    ack_2021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1002_inst_ack_0, ack => convTranspose_CP_34_elements(253)); -- 
    req_2025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(253), ack => WPIPE_Block0_start_1002_inst_req_1); -- 
    -- CP-element group 254:  transition  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (6) 
      -- CP-element group 254: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_update_completed_
      -- CP-element group 254: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_Sample/req
      -- CP-element group 254: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_Update/ack
      -- 
    ack_2026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1002_inst_ack_1, ack => convTranspose_CP_34_elements(254)); -- 
    req_2034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(254), ack => WPIPE_Block0_start_1006_inst_req_0); -- 
    -- CP-element group 255:  transition  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (6) 
      -- CP-element group 255: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_Update/req
      -- CP-element group 255: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_Sample/ack
      -- CP-element group 255: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_update_start_
      -- CP-element group 255: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_sample_completed_
      -- 
    ack_2035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1006_inst_ack_0, ack => convTranspose_CP_34_elements(255)); -- 
    req_2039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(255), ack => WPIPE_Block0_start_1006_inst_req_1); -- 
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_Sample/req
      -- CP-element group 256: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_Update/ack
      -- CP-element group 256: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_update_completed_
      -- 
    ack_2040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1006_inst_ack_1, ack => convTranspose_CP_34_elements(256)); -- 
    req_2048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(256), ack => WPIPE_Block0_start_1010_inst_req_0); -- 
    -- CP-element group 257:  transition  input  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (6) 
      -- CP-element group 257: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_Update/req
      -- CP-element group 257: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_Update/$entry
      -- CP-element group 257: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_Sample/ack
      -- CP-element group 257: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_update_start_
      -- CP-element group 257: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_sample_completed_
      -- 
    ack_2049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1010_inst_ack_0, ack => convTranspose_CP_34_elements(257)); -- 
    req_2053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(257), ack => WPIPE_Block0_start_1010_inst_req_1); -- 
    -- CP-element group 258:  transition  input  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (6) 
      -- CP-element group 258: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_Sample/req
      -- CP-element group 258: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_Update/ack
      -- CP-element group 258: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_update_completed_
      -- 
    ack_2054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1010_inst_ack_1, ack => convTranspose_CP_34_elements(258)); -- 
    req_2062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(258), ack => WPIPE_Block0_start_1013_inst_req_0); -- 
    -- CP-element group 259:  transition  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (6) 
      -- CP-element group 259: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_Update/req
      -- CP-element group 259: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_Sample/ack
      -- CP-element group 259: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_update_start_
      -- CP-element group 259: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_sample_completed_
      -- 
    ack_2063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1013_inst_ack_0, ack => convTranspose_CP_34_elements(259)); -- 
    req_2067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(259), ack => WPIPE_Block0_start_1013_inst_req_1); -- 
    -- CP-element group 260:  transition  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (6) 
      -- CP-element group 260: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_Update/ack
      -- CP-element group 260: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_Sample/req
      -- CP-element group 260: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_update_completed_
      -- 
    ack_2068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1013_inst_ack_1, ack => convTranspose_CP_34_elements(260)); -- 
    req_2076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(260), ack => WPIPE_Block0_start_1016_inst_req_0); -- 
    -- CP-element group 261:  transition  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_update_start_
      -- CP-element group 261: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_sample_completed_
      -- CP-element group 261: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_Sample/ack
      -- CP-element group 261: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_Update/req
      -- 
    ack_2077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1016_inst_ack_0, ack => convTranspose_CP_34_elements(261)); -- 
    req_2081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(261), ack => WPIPE_Block0_start_1016_inst_req_1); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	365 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_Update/ack
      -- CP-element group 262: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_update_completed_
      -- 
    ack_2082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1016_inst_ack_1, ack => convTranspose_CP_34_elements(262)); -- 
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	234 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_update_start_
      -- CP-element group 263: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_Sample/ack
      -- CP-element group 263: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_Update/req
      -- 
    ack_2091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1019_inst_ack_0, ack => convTranspose_CP_34_elements(263)); -- 
    req_2095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(263), ack => WPIPE_Block1_start_1019_inst_req_1); -- 
    -- CP-element group 264:  transition  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (6) 
      -- CP-element group 264: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_Update/ack
      -- CP-element group 264: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_Sample/req
      -- 
    ack_2096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1019_inst_ack_1, ack => convTranspose_CP_34_elements(264)); -- 
    req_2104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(264), ack => WPIPE_Block1_start_1022_inst_req_0); -- 
    -- CP-element group 265:  transition  input  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (6) 
      -- CP-element group 265: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_Update/req
      -- CP-element group 265: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_sample_completed_
      -- CP-element group 265: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_update_start_
      -- CP-element group 265: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_Sample/ack
      -- CP-element group 265: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_Update/$entry
      -- 
    ack_2105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1022_inst_ack_0, ack => convTranspose_CP_34_elements(265)); -- 
    req_2109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(265), ack => WPIPE_Block1_start_1022_inst_req_1); -- 
    -- CP-element group 266:  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (6) 
      -- CP-element group 266: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_Update/ack
      -- CP-element group 266: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_update_completed_
      -- CP-element group 266: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_Sample/req
      -- 
    ack_2110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1022_inst_ack_1, ack => convTranspose_CP_34_elements(266)); -- 
    req_2118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(266), ack => WPIPE_Block1_start_1025_inst_req_0); -- 
    -- CP-element group 267:  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (6) 
      -- CP-element group 267: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_update_start_
      -- CP-element group 267: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_Sample/ack
      -- CP-element group 267: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_Update/req
      -- 
    ack_2119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1025_inst_ack_0, ack => convTranspose_CP_34_elements(267)); -- 
    req_2123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(267), ack => WPIPE_Block1_start_1025_inst_req_1); -- 
    -- CP-element group 268:  transition  input  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (6) 
      -- CP-element group 268: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_update_completed_
      -- CP-element group 268: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_Update/ack
      -- CP-element group 268: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_Sample/req
      -- CP-element group 268: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_Sample/$entry
      -- 
    ack_2124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1025_inst_ack_1, ack => convTranspose_CP_34_elements(268)); -- 
    req_2132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(268), ack => WPIPE_Block1_start_1028_inst_req_0); -- 
    -- CP-element group 269:  transition  input  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (6) 
      -- CP-element group 269: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_Update/req
      -- CP-element group 269: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_Sample/ack
      -- CP-element group 269: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_update_start_
      -- CP-element group 269: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_sample_completed_
      -- 
    ack_2133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1028_inst_ack_0, ack => convTranspose_CP_34_elements(269)); -- 
    req_2137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(269), ack => WPIPE_Block1_start_1028_inst_req_1); -- 
    -- CP-element group 270:  transition  input  output  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (6) 
      -- CP-element group 270: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_Sample/req
      -- CP-element group 270: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_Sample/$entry
      -- CP-element group 270: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_sample_start_
      -- CP-element group 270: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_Update/ack
      -- CP-element group 270: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_update_completed_
      -- 
    ack_2138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1028_inst_ack_1, ack => convTranspose_CP_34_elements(270)); -- 
    req_2146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(270), ack => WPIPE_Block1_start_1031_inst_req_0); -- 
    -- CP-element group 271:  transition  input  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (6) 
      -- CP-element group 271: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_Update/req
      -- CP-element group 271: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_Sample/ack
      -- CP-element group 271: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_update_start_
      -- CP-element group 271: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_sample_completed_
      -- 
    ack_2147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1031_inst_ack_0, ack => convTranspose_CP_34_elements(271)); -- 
    req_2151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(271), ack => WPIPE_Block1_start_1031_inst_req_1); -- 
    -- CP-element group 272:  transition  input  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (6) 
      -- CP-element group 272: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_Update/ack
      -- CP-element group 272: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_Sample/req
      -- CP-element group 272: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_Update/$exit
      -- CP-element group 272: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_update_completed_
      -- 
    ack_2152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1031_inst_ack_1, ack => convTranspose_CP_34_elements(272)); -- 
    req_2160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(272), ack => WPIPE_Block1_start_1034_inst_req_0); -- 
    -- CP-element group 273:  transition  input  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (6) 
      -- CP-element group 273: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_Update/req
      -- CP-element group 273: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_sample_completed_
      -- CP-element group 273: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_update_start_
      -- CP-element group 273: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_Sample/ack
      -- 
    ack_2161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1034_inst_ack_0, ack => convTranspose_CP_34_elements(273)); -- 
    req_2165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(273), ack => WPIPE_Block1_start_1034_inst_req_1); -- 
    -- CP-element group 274:  transition  input  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (6) 
      -- CP-element group 274: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_update_completed_
      -- CP-element group 274: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_Update/ack
      -- CP-element group 274: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_Sample/req
      -- CP-element group 274: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_Sample/$entry
      -- 
    ack_2166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1034_inst_ack_1, ack => convTranspose_CP_34_elements(274)); -- 
    req_2174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(274), ack => WPIPE_Block1_start_1037_inst_req_0); -- 
    -- CP-element group 275:  transition  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (6) 
      -- CP-element group 275: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_sample_completed_
      -- CP-element group 275: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_update_start_
      -- CP-element group 275: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_Update/req
      -- CP-element group 275: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_Sample/ack
      -- CP-element group 275: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_Sample/$exit
      -- 
    ack_2175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1037_inst_ack_0, ack => convTranspose_CP_34_elements(275)); -- 
    req_2179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(275), ack => WPIPE_Block1_start_1037_inst_req_1); -- 
    -- CP-element group 276:  transition  input  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (6) 
      -- CP-element group 276: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_update_completed_
      -- CP-element group 276: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_Sample/req
      -- CP-element group 276: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_Update/ack
      -- CP-element group 276: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_Update/$exit
      -- 
    ack_2180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1037_inst_ack_1, ack => convTranspose_CP_34_elements(276)); -- 
    req_2188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(276), ack => WPIPE_Block1_start_1040_inst_req_0); -- 
    -- CP-element group 277:  transition  input  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (6) 
      -- CP-element group 277: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_Update/req
      -- CP-element group 277: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_Sample/ack
      -- CP-element group 277: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_update_start_
      -- CP-element group 277: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_sample_completed_
      -- 
    ack_2189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1040_inst_ack_0, ack => convTranspose_CP_34_elements(277)); -- 
    req_2193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(277), ack => WPIPE_Block1_start_1040_inst_req_1); -- 
    -- CP-element group 278:  transition  input  output  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (6) 
      -- CP-element group 278: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_Sample/req
      -- CP-element group 278: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_Sample/$entry
      -- CP-element group 278: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_sample_start_
      -- CP-element group 278: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_Update/ack
      -- CP-element group 278: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_update_completed_
      -- 
    ack_2194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1040_inst_ack_1, ack => convTranspose_CP_34_elements(278)); -- 
    req_2202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(278), ack => WPIPE_Block1_start_1043_inst_req_0); -- 
    -- CP-element group 279:  transition  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (6) 
      -- CP-element group 279: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_Update/req
      -- CP-element group 279: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_Sample/ack
      -- CP-element group 279: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_update_start_
      -- CP-element group 279: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_sample_completed_
      -- 
    ack_2203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1043_inst_ack_0, ack => convTranspose_CP_34_elements(279)); -- 
    req_2207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(279), ack => WPIPE_Block1_start_1043_inst_req_1); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	283 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_Update/ack
      -- CP-element group 280: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_update_completed_
      -- 
    ack_2208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1043_inst_ack_1, ack => convTranspose_CP_34_elements(280)); -- 
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	234 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_Sample/ra
      -- CP-element group 281: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_sample_completed_
      -- 
    ra_2217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1054_inst_ack_0, ack => convTranspose_CP_34_elements(281)); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	234 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_Update/ca
      -- CP-element group 282: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_update_completed_
      -- 
    ca_2222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1054_inst_ack_1, ack => convTranspose_CP_34_elements(282)); -- 
    -- CP-element group 283:  join  transition  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	280 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_Sample/req
      -- CP-element group 283: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_sample_start_
      -- 
    req_2230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(283), ack => WPIPE_Block1_start_1056_inst_req_0); -- 
    convTranspose_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(280) & convTranspose_CP_34_elements(282);
      gj_convTranspose_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  transition  input  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (6) 
      -- CP-element group 284: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_Sample/$exit
      -- CP-element group 284: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_Sample/ack
      -- CP-element group 284: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_update_start_
      -- CP-element group 284: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_Update/req
      -- CP-element group 284: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_sample_completed_
      -- 
    ack_2231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1056_inst_ack_0, ack => convTranspose_CP_34_elements(284)); -- 
    req_2235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(284), ack => WPIPE_Block1_start_1056_inst_req_1); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	288 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_update_completed_
      -- CP-element group 285: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_Update/$exit
      -- CP-element group 285: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_Update/ack
      -- 
    ack_2236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1056_inst_ack_1, ack => convTranspose_CP_34_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	234 
    -- CP-element group 286: successors 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_Sample/ra
      -- CP-element group 286: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_Sample/$exit
      -- CP-element group 286: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_sample_completed_
      -- 
    ra_2245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1061_inst_ack_0, ack => convTranspose_CP_34_elements(286)); -- 
    -- CP-element group 287:  transition  input  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	234 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_Update/ca
      -- CP-element group 287: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_Update/$exit
      -- CP-element group 287: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_update_completed_
      -- 
    ca_2250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1061_inst_ack_1, ack => convTranspose_CP_34_elements(287)); -- 
    -- CP-element group 288:  join  transition  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	285 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_Sample/req
      -- CP-element group 288: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_sample_start_
      -- 
    req_2258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(288), ack => WPIPE_Block1_start_1063_inst_req_0); -- 
    convTranspose_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(285) & convTranspose_CP_34_elements(287);
      gj_convTranspose_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  transition  input  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (6) 
      -- CP-element group 289: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_update_start_
      -- CP-element group 289: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_Sample/ack
      -- CP-element group 289: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_Update/req
      -- CP-element group 289: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_sample_completed_
      -- 
    ack_2259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1063_inst_ack_0, ack => convTranspose_CP_34_elements(289)); -- 
    req_2263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(289), ack => WPIPE_Block1_start_1063_inst_req_1); -- 
    -- CP-element group 290:  transition  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (6) 
      -- CP-element group 290: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_update_completed_
      -- CP-element group 290: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_Update/$exit
      -- CP-element group 290: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_Update/ack
      -- CP-element group 290: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_Sample/req
      -- CP-element group 290: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_sample_start_
      -- 
    ack_2264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1063_inst_ack_1, ack => convTranspose_CP_34_elements(290)); -- 
    req_2272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(290), ack => WPIPE_Block1_start_1066_inst_req_0); -- 
    -- CP-element group 291:  transition  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_Update/req
      -- CP-element group 291: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_update_start_
      -- CP-element group 291: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_sample_completed_
      -- 
    ack_2273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1066_inst_ack_0, ack => convTranspose_CP_34_elements(291)); -- 
    req_2277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(291), ack => WPIPE_Block1_start_1066_inst_req_1); -- 
    -- CP-element group 292:  transition  input  output  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (6) 
      -- CP-element group 292: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_Sample/$entry
      -- CP-element group 292: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_Sample/req
      -- CP-element group 292: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_Update/ack
      -- CP-element group 292: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_sample_start_
      -- CP-element group 292: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_update_completed_
      -- 
    ack_2278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1066_inst_ack_1, ack => convTranspose_CP_34_elements(292)); -- 
    req_2286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(292), ack => WPIPE_Block1_start_1069_inst_req_0); -- 
    -- CP-element group 293:  transition  input  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (6) 
      -- CP-element group 293: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_Sample/$exit
      -- CP-element group 293: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_Sample/ack
      -- CP-element group 293: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_update_start_
      -- CP-element group 293: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_sample_completed_
      -- CP-element group 293: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_Update/req
      -- 
    ack_2287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1069_inst_ack_0, ack => convTranspose_CP_34_elements(293)); -- 
    req_2291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(293), ack => WPIPE_Block1_start_1069_inst_req_1); -- 
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_Sample/req
      -- CP-element group 294: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_update_completed_
      -- CP-element group 294: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_sample_start_
      -- CP-element group 294: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_Update/$exit
      -- CP-element group 294: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_Update/ack
      -- 
    ack_2292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1069_inst_ack_1, ack => convTranspose_CP_34_elements(294)); -- 
    req_2300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(294), ack => WPIPE_Block1_start_1072_inst_req_0); -- 
    -- CP-element group 295:  transition  input  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (6) 
      -- CP-element group 295: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_Update/req
      -- CP-element group 295: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_Sample/ack
      -- CP-element group 295: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_update_start_
      -- CP-element group 295: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_sample_completed_
      -- 
    ack_2301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1072_inst_ack_0, ack => convTranspose_CP_34_elements(295)); -- 
    req_2305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(295), ack => WPIPE_Block1_start_1072_inst_req_1); -- 
    -- CP-element group 296:  transition  input  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	365 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_Update/ack
      -- CP-element group 296: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_update_completed_
      -- 
    ack_2306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1072_inst_ack_1, ack => convTranspose_CP_34_elements(296)); -- 
    -- CP-element group 297:  transition  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	234 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (6) 
      -- CP-element group 297: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_Update/req
      -- CP-element group 297: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_Sample/ack
      -- CP-element group 297: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_update_start_
      -- CP-element group 297: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_sample_completed_
      -- 
    ack_2315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1075_inst_ack_0, ack => convTranspose_CP_34_elements(297)); -- 
    req_2319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(297), ack => WPIPE_Block2_start_1075_inst_req_1); -- 
    -- CP-element group 298:  transition  input  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (6) 
      -- CP-element group 298: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_Update/ack
      -- CP-element group 298: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_Sample/req
      -- CP-element group 298: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_update_completed_
      -- CP-element group 298: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_sample_start_
      -- 
    ack_2320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1075_inst_ack_1, ack => convTranspose_CP_34_elements(298)); -- 
    req_2328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(298), ack => WPIPE_Block2_start_1078_inst_req_0); -- 
    -- CP-element group 299:  transition  input  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (6) 
      -- CP-element group 299: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_Update/req
      -- CP-element group 299: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_Sample/ack
      -- CP-element group 299: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_update_start_
      -- CP-element group 299: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_sample_completed_
      -- 
    ack_2329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1078_inst_ack_0, ack => convTranspose_CP_34_elements(299)); -- 
    req_2333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(299), ack => WPIPE_Block2_start_1078_inst_req_1); -- 
    -- CP-element group 300:  transition  input  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (6) 
      -- CP-element group 300: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_Update/ack
      -- CP-element group 300: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_Sample/req
      -- CP-element group 300: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_Sample/$entry
      -- CP-element group 300: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_update_completed_
      -- CP-element group 300: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_sample_start_
      -- 
    ack_2334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1078_inst_ack_1, ack => convTranspose_CP_34_elements(300)); -- 
    req_2342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(300), ack => WPIPE_Block2_start_1081_inst_req_0); -- 
    -- CP-element group 301:  transition  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (6) 
      -- CP-element group 301: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_Update/req
      -- CP-element group 301: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_Sample/ack
      -- CP-element group 301: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_Sample/$exit
      -- CP-element group 301: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_update_start_
      -- CP-element group 301: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_sample_completed_
      -- 
    ack_2343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1081_inst_ack_0, ack => convTranspose_CP_34_elements(301)); -- 
    req_2347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(301), ack => WPIPE_Block2_start_1081_inst_req_1); -- 
    -- CP-element group 302:  transition  input  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (6) 
      -- CP-element group 302: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_Update/ack
      -- CP-element group 302: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_Sample/req
      -- CP-element group 302: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_Update/$exit
      -- CP-element group 302: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_update_completed_
      -- 
    ack_2348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1081_inst_ack_1, ack => convTranspose_CP_34_elements(302)); -- 
    req_2356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(302), ack => WPIPE_Block2_start_1084_inst_req_0); -- 
    -- CP-element group 303:  transition  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_Update/req
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_update_start_
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_sample_completed_
      -- 
    ack_2357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1084_inst_ack_0, ack => convTranspose_CP_34_elements(303)); -- 
    req_2361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(303), ack => WPIPE_Block2_start_1084_inst_req_1); -- 
    -- CP-element group 304:  transition  input  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (6) 
      -- CP-element group 304: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_Update/ack
      -- CP-element group 304: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_sample_start_
      -- CP-element group 304: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_Sample/req
      -- CP-element group 304: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_Sample/$entry
      -- 
    ack_2362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1084_inst_ack_1, ack => convTranspose_CP_34_elements(304)); -- 
    req_2370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(304), ack => WPIPE_Block2_start_1087_inst_req_0); -- 
    -- CP-element group 305:  transition  input  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (6) 
      -- CP-element group 305: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_update_start_
      -- CP-element group 305: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_Update/req
      -- CP-element group 305: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_sample_completed_
      -- CP-element group 305: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_Update/$entry
      -- CP-element group 305: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_Sample/ack
      -- CP-element group 305: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_Sample/$exit
      -- 
    ack_2371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1087_inst_ack_0, ack => convTranspose_CP_34_elements(305)); -- 
    req_2375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(305), ack => WPIPE_Block2_start_1087_inst_req_1); -- 
    -- CP-element group 306:  transition  input  output  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (6) 
      -- CP-element group 306: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_Update/ack
      -- CP-element group 306: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_Sample/req
      -- CP-element group 306: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_Sample/$entry
      -- CP-element group 306: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_Update/$exit
      -- CP-element group 306: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_sample_start_
      -- CP-element group 306: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_update_completed_
      -- 
    ack_2376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1087_inst_ack_1, ack => convTranspose_CP_34_elements(306)); -- 
    req_2384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(306), ack => WPIPE_Block2_start_1090_inst_req_0); -- 
    -- CP-element group 307:  transition  input  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (6) 
      -- CP-element group 307: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_Sample/ack
      -- CP-element group 307: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_update_start_
      -- CP-element group 307: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_sample_completed_
      -- CP-element group 307: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_Update/req
      -- CP-element group 307: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_Update/$entry
      -- 
    ack_2385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1090_inst_ack_0, ack => convTranspose_CP_34_elements(307)); -- 
    req_2389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(307), ack => WPIPE_Block2_start_1090_inst_req_1); -- 
    -- CP-element group 308:  transition  input  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (6) 
      -- CP-element group 308: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_Update/ack
      -- CP-element group 308: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_Sample/req
      -- 
    ack_2390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1090_inst_ack_1, ack => convTranspose_CP_34_elements(308)); -- 
    req_2398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(308), ack => WPIPE_Block2_start_1093_inst_req_0); -- 
    -- CP-element group 309:  transition  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (6) 
      -- CP-element group 309: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_update_start_
      -- CP-element group 309: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_sample_completed_
      -- CP-element group 309: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_Sample/$exit
      -- CP-element group 309: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_Sample/ack
      -- CP-element group 309: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_Update/req
      -- 
    ack_2399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1093_inst_ack_0, ack => convTranspose_CP_34_elements(309)); -- 
    req_2403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(309), ack => WPIPE_Block2_start_1093_inst_req_1); -- 
    -- CP-element group 310:  transition  input  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (6) 
      -- CP-element group 310: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_update_completed_
      -- CP-element group 310: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_Update/$exit
      -- CP-element group 310: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_Update/ack
      -- CP-element group 310: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_sample_start_
      -- CP-element group 310: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_Sample/req
      -- 
    ack_2404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1093_inst_ack_1, ack => convTranspose_CP_34_elements(310)); -- 
    req_2412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(310), ack => WPIPE_Block2_start_1096_inst_req_0); -- 
    -- CP-element group 311:  transition  input  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (6) 
      -- CP-element group 311: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_sample_completed_
      -- CP-element group 311: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_update_start_
      -- CP-element group 311: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_Sample/ack
      -- CP-element group 311: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_Update/req
      -- 
    ack_2413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1096_inst_ack_0, ack => convTranspose_CP_34_elements(311)); -- 
    req_2417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(311), ack => WPIPE_Block2_start_1096_inst_req_1); -- 
    -- CP-element group 312:  transition  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (6) 
      -- CP-element group 312: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_Update/ack
      -- CP-element group 312: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_sample_start_
      -- CP-element group 312: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_Sample/$entry
      -- CP-element group 312: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_Sample/req
      -- 
    ack_2418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1096_inst_ack_1, ack => convTranspose_CP_34_elements(312)); -- 
    req_2426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(312), ack => WPIPE_Block2_start_1099_inst_req_0); -- 
    -- CP-element group 313:  transition  input  output  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (6) 
      -- CP-element group 313: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_sample_completed_
      -- CP-element group 313: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_update_start_
      -- CP-element group 313: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_Sample/$exit
      -- CP-element group 313: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_Sample/ack
      -- CP-element group 313: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_Update/$entry
      -- CP-element group 313: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_Update/req
      -- 
    ack_2427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1099_inst_ack_0, ack => convTranspose_CP_34_elements(313)); -- 
    req_2431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(313), ack => WPIPE_Block2_start_1099_inst_req_1); -- 
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	317 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_update_completed_
      -- CP-element group 314: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_Update/$exit
      -- CP-element group 314: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_Update/ack
      -- 
    ack_2432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1099_inst_ack_1, ack => convTranspose_CP_34_elements(314)); -- 
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	234 
    -- CP-element group 315: successors 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_Sample/ra
      -- 
    ra_2441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1110_inst_ack_0, ack => convTranspose_CP_34_elements(315)); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	234 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_Update/ca
      -- 
    ca_2446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1110_inst_ack_1, ack => convTranspose_CP_34_elements(316)); -- 
    -- CP-element group 317:  join  transition  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	314 
    -- CP-element group 317: 	316 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_Sample/req
      -- 
    req_2454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(317), ack => WPIPE_Block2_start_1112_inst_req_0); -- 
    convTranspose_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(314) & convTranspose_CP_34_elements(316);
      gj_convTranspose_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  transition  input  output  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (6) 
      -- CP-element group 318: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_sample_completed_
      -- CP-element group 318: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_update_start_
      -- CP-element group 318: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_Sample/$exit
      -- CP-element group 318: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_Sample/ack
      -- CP-element group 318: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_Update/$entry
      -- CP-element group 318: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_Update/req
      -- 
    ack_2455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1112_inst_ack_0, ack => convTranspose_CP_34_elements(318)); -- 
    req_2459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(318), ack => WPIPE_Block2_start_1112_inst_req_1); -- 
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	322 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_update_completed_
      -- CP-element group 319: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_Update/$exit
      -- CP-element group 319: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_Update/ack
      -- 
    ack_2460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1112_inst_ack_1, ack => convTranspose_CP_34_elements(319)); -- 
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	234 
    -- CP-element group 320: successors 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_sample_completed_
      -- CP-element group 320: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_Sample/ra
      -- 
    ra_2469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1117_inst_ack_0, ack => convTranspose_CP_34_elements(320)); -- 
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	234 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_update_completed_
      -- CP-element group 321: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_Update/ca
      -- 
    ca_2474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1117_inst_ack_1, ack => convTranspose_CP_34_elements(321)); -- 
    -- CP-element group 322:  join  transition  output  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	319 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_sample_start_
      -- CP-element group 322: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_Sample/req
      -- 
    req_2482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(322), ack => WPIPE_Block2_start_1119_inst_req_0); -- 
    convTranspose_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(319) & convTranspose_CP_34_elements(321);
      gj_convTranspose_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  transition  input  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (6) 
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_sample_completed_
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_update_start_
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_Sample/ack
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_Update/req
      -- 
    ack_2483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1119_inst_ack_0, ack => convTranspose_CP_34_elements(323)); -- 
    req_2487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(323), ack => WPIPE_Block2_start_1119_inst_req_1); -- 
    -- CP-element group 324:  transition  input  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (6) 
      -- CP-element group 324: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_update_completed_
      -- CP-element group 324: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_Update/ack
      -- CP-element group 324: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_sample_start_
      -- CP-element group 324: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_Sample/$entry
      -- CP-element group 324: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_Sample/req
      -- 
    ack_2488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1119_inst_ack_1, ack => convTranspose_CP_34_elements(324)); -- 
    req_2496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(324), ack => WPIPE_Block2_start_1122_inst_req_0); -- 
    -- CP-element group 325:  transition  input  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (6) 
      -- CP-element group 325: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_sample_completed_
      -- CP-element group 325: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_update_start_
      -- CP-element group 325: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_Sample/$exit
      -- CP-element group 325: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_Sample/ack
      -- CP-element group 325: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_Update/req
      -- 
    ack_2497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1122_inst_ack_0, ack => convTranspose_CP_34_elements(325)); -- 
    req_2501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(325), ack => WPIPE_Block2_start_1122_inst_req_1); -- 
    -- CP-element group 326:  transition  input  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (6) 
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_update_completed_
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_Update/$exit
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_Update/ack
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_Sample/req
      -- 
    ack_2502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1122_inst_ack_1, ack => convTranspose_CP_34_elements(326)); -- 
    req_2510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(326), ack => WPIPE_Block2_start_1125_inst_req_0); -- 
    -- CP-element group 327:  transition  input  output  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (6) 
      -- CP-element group 327: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_update_start_
      -- CP-element group 327: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_Sample/ack
      -- CP-element group 327: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_Update/$entry
      -- CP-element group 327: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_Update/req
      -- 
    ack_2511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1125_inst_ack_0, ack => convTranspose_CP_34_elements(327)); -- 
    req_2515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(327), ack => WPIPE_Block2_start_1125_inst_req_1); -- 
    -- CP-element group 328:  transition  input  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328:  members (6) 
      -- CP-element group 328: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_Update/ack
      -- CP-element group 328: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_sample_start_
      -- CP-element group 328: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_Sample/$entry
      -- CP-element group 328: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_Sample/req
      -- 
    ack_2516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1125_inst_ack_1, ack => convTranspose_CP_34_elements(328)); -- 
    req_2524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(328), ack => WPIPE_Block2_start_1128_inst_req_0); -- 
    -- CP-element group 329:  transition  input  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	330 
    -- CP-element group 329:  members (6) 
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_sample_completed_
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_update_start_
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_Sample/$exit
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_Sample/ack
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_Update/req
      -- 
    ack_2525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1128_inst_ack_0, ack => convTranspose_CP_34_elements(329)); -- 
    req_2529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(329), ack => WPIPE_Block2_start_1128_inst_req_1); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	329 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	365 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_update_completed_
      -- CP-element group 330: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_Update/$exit
      -- CP-element group 330: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_Update/ack
      -- 
    ack_2530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1128_inst_ack_1, ack => convTranspose_CP_34_elements(330)); -- 
    -- CP-element group 331:  transition  input  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	234 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (6) 
      -- CP-element group 331: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_sample_completed_
      -- CP-element group 331: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_update_start_
      -- CP-element group 331: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_Sample/ack
      -- CP-element group 331: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_Update/$entry
      -- CP-element group 331: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_Update/req
      -- 
    ack_2539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1131_inst_ack_0, ack => convTranspose_CP_34_elements(331)); -- 
    req_2543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(331), ack => WPIPE_Block3_start_1131_inst_req_1); -- 
    -- CP-element group 332:  transition  input  output  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (6) 
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_update_completed_
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_Update/ack
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_sample_start_
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_Sample/$entry
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_Sample/req
      -- 
    ack_2544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1131_inst_ack_1, ack => convTranspose_CP_34_elements(332)); -- 
    req_2552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(332), ack => WPIPE_Block3_start_1134_inst_req_0); -- 
    -- CP-element group 333:  transition  input  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (6) 
      -- CP-element group 333: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_sample_completed_
      -- CP-element group 333: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_update_start_
      -- CP-element group 333: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_Sample/$exit
      -- CP-element group 333: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_Sample/ack
      -- CP-element group 333: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_Update/req
      -- 
    ack_2553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1134_inst_ack_0, ack => convTranspose_CP_34_elements(333)); -- 
    req_2557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(333), ack => WPIPE_Block3_start_1134_inst_req_1); -- 
    -- CP-element group 334:  transition  input  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (6) 
      -- CP-element group 334: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_update_completed_
      -- CP-element group 334: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_Update/$exit
      -- CP-element group 334: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_Update/ack
      -- CP-element group 334: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_sample_start_
      -- CP-element group 334: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_Sample/$entry
      -- CP-element group 334: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_Sample/req
      -- 
    ack_2558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1134_inst_ack_1, ack => convTranspose_CP_34_elements(334)); -- 
    req_2566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(334), ack => WPIPE_Block3_start_1137_inst_req_0); -- 
    -- CP-element group 335:  transition  input  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (6) 
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_sample_completed_
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_update_start_
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_Sample/ack
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_Update/req
      -- 
    ack_2567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1137_inst_ack_0, ack => convTranspose_CP_34_elements(335)); -- 
    req_2571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(335), ack => WPIPE_Block3_start_1137_inst_req_1); -- 
    -- CP-element group 336:  transition  input  output  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336:  members (6) 
      -- CP-element group 336: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_update_completed_
      -- CP-element group 336: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_Update/$exit
      -- CP-element group 336: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_Update/ack
      -- CP-element group 336: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_Sample/req
      -- 
    ack_2572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1137_inst_ack_1, ack => convTranspose_CP_34_elements(336)); -- 
    req_2580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(336), ack => WPIPE_Block3_start_1140_inst_req_0); -- 
    -- CP-element group 337:  transition  input  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (6) 
      -- CP-element group 337: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_sample_completed_
      -- CP-element group 337: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_update_start_
      -- CP-element group 337: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_Sample/$exit
      -- CP-element group 337: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_Sample/ack
      -- CP-element group 337: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_Update/req
      -- 
    ack_2581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1140_inst_ack_0, ack => convTranspose_CP_34_elements(337)); -- 
    req_2585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(337), ack => WPIPE_Block3_start_1140_inst_req_1); -- 
    -- CP-element group 338:  transition  input  output  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	337 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338:  members (6) 
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_update_completed_
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_Update/ack
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_sample_start_
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_Sample/$entry
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_Sample/req
      -- 
    ack_2586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1140_inst_ack_1, ack => convTranspose_CP_34_elements(338)); -- 
    req_2594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(338), ack => WPIPE_Block3_start_1143_inst_req_0); -- 
    -- CP-element group 339:  transition  input  output  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	338 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339:  members (6) 
      -- CP-element group 339: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_sample_completed_
      -- CP-element group 339: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_update_start_
      -- CP-element group 339: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_Sample/$exit
      -- CP-element group 339: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_Sample/ack
      -- CP-element group 339: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_Update/req
      -- 
    ack_2595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1143_inst_ack_0, ack => convTranspose_CP_34_elements(339)); -- 
    req_2599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(339), ack => WPIPE_Block3_start_1143_inst_req_1); -- 
    -- CP-element group 340:  transition  input  output  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (6) 
      -- CP-element group 340: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_update_completed_
      -- CP-element group 340: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_Update/$exit
      -- CP-element group 340: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_Update/ack
      -- CP-element group 340: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_sample_start_
      -- CP-element group 340: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_Sample/$entry
      -- CP-element group 340: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_Sample/req
      -- 
    ack_2600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1143_inst_ack_1, ack => convTranspose_CP_34_elements(340)); -- 
    req_2608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(340), ack => WPIPE_Block3_start_1146_inst_req_0); -- 
    -- CP-element group 341:  transition  input  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (6) 
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_sample_completed_
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_update_start_
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_Sample/$exit
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_Sample/ack
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_Update/req
      -- 
    ack_2609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1146_inst_ack_0, ack => convTranspose_CP_34_elements(341)); -- 
    req_2613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(341), ack => WPIPE_Block3_start_1146_inst_req_1); -- 
    -- CP-element group 342:  transition  input  output  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	343 
    -- CP-element group 342:  members (6) 
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_update_completed_
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_Update/$exit
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_Update/ack
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_sample_start_
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_Sample/req
      -- 
    ack_2614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1146_inst_ack_1, ack => convTranspose_CP_34_elements(342)); -- 
    req_2622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(342), ack => WPIPE_Block3_start_1149_inst_req_0); -- 
    -- CP-element group 343:  transition  input  output  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	342 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343:  members (6) 
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_sample_completed_
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_update_start_
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_Sample/$exit
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_Sample/ack
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_Update/req
      -- 
    ack_2623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1149_inst_ack_0, ack => convTranspose_CP_34_elements(343)); -- 
    req_2627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(343), ack => WPIPE_Block3_start_1149_inst_req_1); -- 
    -- CP-element group 344:  transition  input  output  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	343 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	345 
    -- CP-element group 344:  members (6) 
      -- CP-element group 344: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_Update/$exit
      -- CP-element group 344: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_Update/ack
      -- CP-element group 344: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_sample_start_
      -- CP-element group 344: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_Sample/$entry
      -- CP-element group 344: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_Sample/req
      -- 
    ack_2628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1149_inst_ack_1, ack => convTranspose_CP_34_elements(344)); -- 
    req_2636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(344), ack => WPIPE_Block3_start_1152_inst_req_0); -- 
    -- CP-element group 345:  transition  input  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	344 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345:  members (6) 
      -- CP-element group 345: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_sample_completed_
      -- CP-element group 345: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_update_start_
      -- CP-element group 345: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_Sample/$exit
      -- CP-element group 345: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_Sample/ack
      -- CP-element group 345: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_Update/req
      -- 
    ack_2637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1152_inst_ack_0, ack => convTranspose_CP_34_elements(345)); -- 
    req_2641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(345), ack => WPIPE_Block3_start_1152_inst_req_1); -- 
    -- CP-element group 346:  transition  input  output  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	347 
    -- CP-element group 346:  members (6) 
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_update_completed_
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_Update/$exit
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_Update/ack
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_sample_start_
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_Sample/$entry
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_Sample/req
      -- 
    ack_2642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1152_inst_ack_1, ack => convTranspose_CP_34_elements(346)); -- 
    req_2650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(346), ack => WPIPE_Block3_start_1155_inst_req_0); -- 
    -- CP-element group 347:  transition  input  output  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	346 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (6) 
      -- CP-element group 347: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_sample_completed_
      -- CP-element group 347: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_update_start_
      -- CP-element group 347: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_Sample/$exit
      -- CP-element group 347: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_Sample/ack
      -- CP-element group 347: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_Update/$entry
      -- CP-element group 347: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_Update/req
      -- 
    ack_2651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1155_inst_ack_0, ack => convTranspose_CP_34_elements(347)); -- 
    req_2655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(347), ack => WPIPE_Block3_start_1155_inst_req_1); -- 
    -- CP-element group 348:  transition  input  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	351 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_update_completed_
      -- CP-element group 348: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_Update/ack
      -- 
    ack_2656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1155_inst_ack_1, ack => convTranspose_CP_34_elements(348)); -- 
    -- CP-element group 349:  transition  input  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	234 
    -- CP-element group 349: successors 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_sample_completed_
      -- CP-element group 349: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_Sample/$exit
      -- CP-element group 349: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_Sample/ra
      -- 
    ra_2665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1166_inst_ack_0, ack => convTranspose_CP_34_elements(349)); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	234 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	351 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_update_completed_
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_Update/$exit
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_Update/ca
      -- 
    ca_2670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1166_inst_ack_1, ack => convTranspose_CP_34_elements(350)); -- 
    -- CP-element group 351:  join  transition  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	350 
    -- CP-element group 351: 	348 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_sample_start_
      -- CP-element group 351: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_Sample/$entry
      -- CP-element group 351: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_Sample/req
      -- 
    req_2678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(351), ack => WPIPE_Block3_start_1168_inst_req_0); -- 
    convTranspose_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(350) & convTranspose_CP_34_elements(348);
      gj_convTranspose_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  transition  input  output  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (6) 
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_sample_completed_
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_update_start_
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_Sample/ack
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_Update/req
      -- 
    ack_2679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1168_inst_ack_0, ack => convTranspose_CP_34_elements(352)); -- 
    req_2683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(352), ack => WPIPE_Block3_start_1168_inst_req_1); -- 
    -- CP-element group 353:  transition  input  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	356 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_update_completed_
      -- CP-element group 353: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_Update/$exit
      -- CP-element group 353: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_Update/ack
      -- 
    ack_2684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1168_inst_ack_1, ack => convTranspose_CP_34_elements(353)); -- 
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	234 
    -- CP-element group 354: successors 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_sample_completed_
      -- CP-element group 354: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_Sample/$exit
      -- CP-element group 354: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_Sample/ra
      -- 
    ra_2693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1173_inst_ack_0, ack => convTranspose_CP_34_elements(354)); -- 
    -- CP-element group 355:  transition  input  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	234 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_update_completed_
      -- CP-element group 355: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_Update/$exit
      -- CP-element group 355: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_Update/ca
      -- 
    ca_2698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1173_inst_ack_1, ack => convTranspose_CP_34_elements(355)); -- 
    -- CP-element group 356:  join  transition  output  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	353 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	357 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_sample_start_
      -- CP-element group 356: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_Sample/$entry
      -- CP-element group 356: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_Sample/req
      -- 
    req_2706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(356), ack => WPIPE_Block3_start_1175_inst_req_0); -- 
    convTranspose_cp_element_group_356: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_356"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(353) & convTranspose_CP_34_elements(355);
      gj_convTranspose_cp_element_group_356 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(356), clk => clk, reset => reset); --
    end block;
    -- CP-element group 357:  transition  input  output  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	356 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (6) 
      -- CP-element group 357: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_sample_completed_
      -- CP-element group 357: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_update_start_
      -- CP-element group 357: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_Sample/$exit
      -- CP-element group 357: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_Sample/ack
      -- CP-element group 357: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_Update/$entry
      -- CP-element group 357: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_Update/req
      -- 
    ack_2707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1175_inst_ack_0, ack => convTranspose_CP_34_elements(357)); -- 
    req_2711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(357), ack => WPIPE_Block3_start_1175_inst_req_1); -- 
    -- CP-element group 358:  transition  input  output  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (6) 
      -- CP-element group 358: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_update_completed_
      -- CP-element group 358: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_Update/$exit
      -- CP-element group 358: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_Update/ack
      -- CP-element group 358: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_sample_start_
      -- CP-element group 358: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_Sample/$entry
      -- CP-element group 358: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_Sample/req
      -- 
    ack_2712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1175_inst_ack_1, ack => convTranspose_CP_34_elements(358)); -- 
    req_2720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(358), ack => WPIPE_Block3_start_1178_inst_req_0); -- 
    -- CP-element group 359:  transition  input  output  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	360 
    -- CP-element group 359:  members (6) 
      -- CP-element group 359: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_sample_completed_
      -- CP-element group 359: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_update_start_
      -- CP-element group 359: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_Sample/$exit
      -- CP-element group 359: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_Sample/ack
      -- CP-element group 359: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_Update/req
      -- 
    ack_2721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1178_inst_ack_0, ack => convTranspose_CP_34_elements(359)); -- 
    req_2725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(359), ack => WPIPE_Block3_start_1178_inst_req_1); -- 
    -- CP-element group 360:  transition  input  output  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	359 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360:  members (6) 
      -- CP-element group 360: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_update_completed_
      -- CP-element group 360: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_Update/$exit
      -- CP-element group 360: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_Update/ack
      -- CP-element group 360: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_sample_start_
      -- CP-element group 360: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_Sample/$entry
      -- CP-element group 360: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_Sample/req
      -- 
    ack_2726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1178_inst_ack_1, ack => convTranspose_CP_34_elements(360)); -- 
    req_2734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(360), ack => WPIPE_Block3_start_1181_inst_req_0); -- 
    -- CP-element group 361:  transition  input  output  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	360 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (6) 
      -- CP-element group 361: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_sample_completed_
      -- CP-element group 361: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_update_start_
      -- CP-element group 361: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_Sample/$exit
      -- CP-element group 361: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_Sample/ack
      -- CP-element group 361: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_Update/$entry
      -- CP-element group 361: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_Update/req
      -- 
    ack_2735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1181_inst_ack_0, ack => convTranspose_CP_34_elements(361)); -- 
    req_2739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(361), ack => WPIPE_Block3_start_1181_inst_req_1); -- 
    -- CP-element group 362:  transition  input  output  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362:  members (6) 
      -- CP-element group 362: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_update_completed_
      -- CP-element group 362: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_Update/$exit
      -- CP-element group 362: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_Update/ack
      -- CP-element group 362: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_sample_start_
      -- CP-element group 362: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_Sample/$entry
      -- CP-element group 362: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_Sample/req
      -- 
    ack_2740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1181_inst_ack_1, ack => convTranspose_CP_34_elements(362)); -- 
    req_2748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(362), ack => WPIPE_Block3_start_1184_inst_req_0); -- 
    -- CP-element group 363:  transition  input  output  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (6) 
      -- CP-element group 363: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_sample_completed_
      -- CP-element group 363: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_update_start_
      -- CP-element group 363: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_Sample/$exit
      -- CP-element group 363: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_Sample/ack
      -- CP-element group 363: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_Update/req
      -- 
    ack_2749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1184_inst_ack_0, ack => convTranspose_CP_34_elements(363)); -- 
    req_2753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(363), ack => WPIPE_Block3_start_1184_inst_req_1); -- 
    -- CP-element group 364:  transition  input  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	365 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_update_completed_
      -- CP-element group 364: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_Update/$exit
      -- CP-element group 364: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_Update/ack
      -- 
    ack_2754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1184_inst_ack_1, ack => convTranspose_CP_34_elements(364)); -- 
    -- CP-element group 365:  join  fork  transition  place  output  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	364 
    -- CP-element group 365: 	262 
    -- CP-element group 365: 	296 
    -- CP-element group 365: 	330 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	368 
    -- CP-element group 365: 	370 
    -- CP-element group 365: 	372 
    -- CP-element group 365: 	366 
    -- CP-element group 365:  members (16) 
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186__exit__
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199__entry__
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/$exit
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/$entry
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_sample_start_
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_Sample/rr
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_sample_start_
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_Sample/rr
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_sample_start_
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_Sample/rr
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_sample_start_
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_Sample/rr
      -- 
    rr_2765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(365), ack => RPIPE_Block0_done_1189_inst_req_0); -- 
    rr_2779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(365), ack => RPIPE_Block1_done_1192_inst_req_0); -- 
    rr_2793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(365), ack => RPIPE_Block2_done_1195_inst_req_0); -- 
    rr_2807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(365), ack => RPIPE_Block3_done_1198_inst_req_0); -- 
    convTranspose_cp_element_group_365: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_365"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(364) & convTranspose_CP_34_elements(262) & convTranspose_CP_34_elements(296) & convTranspose_CP_34_elements(330);
      gj_convTranspose_cp_element_group_365 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(365), clk => clk, reset => reset); --
    end block;
    -- CP-element group 366:  transition  input  output  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	367 
    -- CP-element group 366:  members (6) 
      -- CP-element group 366: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_sample_completed_
      -- CP-element group 366: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_update_start_
      -- CP-element group 366: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_Sample/$exit
      -- CP-element group 366: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_Sample/ra
      -- CP-element group 366: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_Update/cr
      -- 
    ra_2766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1189_inst_ack_0, ack => convTranspose_CP_34_elements(366)); -- 
    cr_2770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(366), ack => RPIPE_Block0_done_1189_inst_req_1); -- 
    -- CP-element group 367:  transition  input  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	366 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	374 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_update_completed_
      -- CP-element group 367: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_Update/$exit
      -- CP-element group 367: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_Update/ca
      -- 
    ca_2771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1189_inst_ack_1, ack => convTranspose_CP_34_elements(367)); -- 
    -- CP-element group 368:  transition  input  output  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	365 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	369 
    -- CP-element group 368:  members (6) 
      -- CP-element group 368: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_sample_completed_
      -- CP-element group 368: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_update_start_
      -- CP-element group 368: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_Sample/$exit
      -- CP-element group 368: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_Sample/ra
      -- CP-element group 368: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_Update/cr
      -- 
    ra_2780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1192_inst_ack_0, ack => convTranspose_CP_34_elements(368)); -- 
    cr_2784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(368), ack => RPIPE_Block1_done_1192_inst_req_1); -- 
    -- CP-element group 369:  transition  input  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	368 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	374 
    -- CP-element group 369:  members (3) 
      -- CP-element group 369: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_update_completed_
      -- CP-element group 369: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_Update/$exit
      -- CP-element group 369: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_Update/ca
      -- 
    ca_2785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1192_inst_ack_1, ack => convTranspose_CP_34_elements(369)); -- 
    -- CP-element group 370:  transition  input  output  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	365 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	371 
    -- CP-element group 370:  members (6) 
      -- CP-element group 370: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_sample_completed_
      -- CP-element group 370: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_update_start_
      -- CP-element group 370: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_Sample/$exit
      -- CP-element group 370: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_Sample/ra
      -- CP-element group 370: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_Update/cr
      -- 
    ra_2794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1195_inst_ack_0, ack => convTranspose_CP_34_elements(370)); -- 
    cr_2798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(370), ack => RPIPE_Block2_done_1195_inst_req_1); -- 
    -- CP-element group 371:  transition  input  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	370 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	374 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_update_completed_
      -- CP-element group 371: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_Update/$exit
      -- CP-element group 371: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_Update/ca
      -- 
    ca_2799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1195_inst_ack_1, ack => convTranspose_CP_34_elements(371)); -- 
    -- CP-element group 372:  transition  input  output  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	365 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (6) 
      -- CP-element group 372: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_sample_completed_
      -- CP-element group 372: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_update_start_
      -- CP-element group 372: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_Sample/$exit
      -- CP-element group 372: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_Sample/ra
      -- CP-element group 372: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_Update/cr
      -- 
    ra_2808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1198_inst_ack_0, ack => convTranspose_CP_34_elements(372)); -- 
    cr_2812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(372), ack => RPIPE_Block3_done_1198_inst_req_1); -- 
    -- CP-element group 373:  transition  input  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (3) 
      -- CP-element group 373: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_update_completed_
      -- CP-element group 373: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_Update/$exit
      -- CP-element group 373: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_Update/ca
      -- 
    ca_2813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1198_inst_ack_1, ack => convTranspose_CP_34_elements(373)); -- 
    -- CP-element group 374:  join  fork  transition  place  output  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	367 
    -- CP-element group 374: 	369 
    -- CP-element group 374: 	371 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	375 
    -- CP-element group 374: 	376 
    -- CP-element group 374: 	378 
    -- CP-element group 374: 	380 
    -- CP-element group 374: 	382 
    -- CP-element group 374: 	384 
    -- CP-element group 374: 	386 
    -- CP-element group 374: 	388 
    -- CP-element group 374: 	390 
    -- CP-element group 374: 	392 
    -- CP-element group 374: 	394 
    -- CP-element group 374:  members (37) 
      -- CP-element group 374: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199__exit__
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310__entry__
      -- CP-element group 374: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/$exit
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_sample_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_update_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_Sample/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_Sample/crr
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_Update/ccr
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_update_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_update_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_update_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_update_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_update_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_update_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_update_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_update_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_update_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_Update/cr
      -- 
    crr_2824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => call_stmt_1202_call_req_0); -- 
    ccr_2829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => call_stmt_1202_call_req_1); -- 
    cr_2843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1206_inst_req_1); -- 
    cr_2857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1215_inst_req_1); -- 
    cr_2871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1225_inst_req_1); -- 
    cr_2885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1235_inst_req_1); -- 
    cr_2899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1245_inst_req_1); -- 
    cr_2913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1255_inst_req_1); -- 
    cr_2927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1265_inst_req_1); -- 
    cr_2941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1275_inst_req_1); -- 
    cr_2955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1285_inst_req_1); -- 
    convTranspose_cp_element_group_374: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_374"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(367) & convTranspose_CP_34_elements(369) & convTranspose_CP_34_elements(371) & convTranspose_CP_34_elements(373);
      gj_convTranspose_cp_element_group_374 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(374), clk => clk, reset => reset); --
    end block;
    -- CP-element group 375:  transition  input  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	374 
    -- CP-element group 375: successors 
    -- CP-element group 375:  members (3) 
      -- CP-element group 375: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_sample_completed_
      -- CP-element group 375: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_Sample/$exit
      -- CP-element group 375: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_Sample/cra
      -- 
    cra_2825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1202_call_ack_0, ack => convTranspose_CP_34_elements(375)); -- 
    -- CP-element group 376:  transition  input  output  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	374 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	377 
    -- CP-element group 376:  members (6) 
      -- CP-element group 376: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_update_completed_
      -- CP-element group 376: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_Update/$exit
      -- CP-element group 376: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_Update/cca
      -- CP-element group 376: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_sample_start_
      -- CP-element group 376: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_Sample/$entry
      -- CP-element group 376: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_Sample/rr
      -- 
    cca_2830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1202_call_ack_1, ack => convTranspose_CP_34_elements(376)); -- 
    rr_2838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(376), ack => type_cast_1206_inst_req_0); -- 
    -- CP-element group 377:  transition  input  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	376 
    -- CP-element group 377: successors 
    -- CP-element group 377:  members (3) 
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_sample_completed_
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_Sample/$exit
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_Sample/ra
      -- 
    ra_2839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1206_inst_ack_0, ack => convTranspose_CP_34_elements(377)); -- 
    -- CP-element group 378:  fork  transition  input  output  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	374 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	379 
    -- CP-element group 378: 	381 
    -- CP-element group 378: 	383 
    -- CP-element group 378: 	385 
    -- CP-element group 378: 	387 
    -- CP-element group 378: 	389 
    -- CP-element group 378: 	391 
    -- CP-element group 378: 	393 
    -- CP-element group 378:  members (27) 
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_update_completed_
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_Update/$exit
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_Update/ca
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_Sample/rr
      -- 
    ca_2844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1206_inst_ack_1, ack => convTranspose_CP_34_elements(378)); -- 
    rr_2852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1215_inst_req_0); -- 
    rr_2866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1225_inst_req_0); -- 
    rr_2880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1235_inst_req_0); -- 
    rr_2894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1245_inst_req_0); -- 
    rr_2908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1255_inst_req_0); -- 
    rr_2922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1265_inst_req_0); -- 
    rr_2936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1275_inst_req_0); -- 
    rr_2950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1285_inst_req_0); -- 
    -- CP-element group 379:  transition  input  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	378 
    -- CP-element group 379: successors 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_sample_completed_
      -- CP-element group 379: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_Sample/$exit
      -- CP-element group 379: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_Sample/ra
      -- 
    ra_2853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1215_inst_ack_0, ack => convTranspose_CP_34_elements(379)); -- 
    -- CP-element group 380:  transition  input  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	374 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	415 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_update_completed_
      -- CP-element group 380: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_Update/$exit
      -- CP-element group 380: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_Update/ca
      -- 
    ca_2858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1215_inst_ack_1, ack => convTranspose_CP_34_elements(380)); -- 
    -- CP-element group 381:  transition  input  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	378 
    -- CP-element group 381: successors 
    -- CP-element group 381:  members (3) 
      -- CP-element group 381: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_sample_completed_
      -- CP-element group 381: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_Sample/$exit
      -- CP-element group 381: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_Sample/ra
      -- 
    ra_2867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1225_inst_ack_0, ack => convTranspose_CP_34_elements(381)); -- 
    -- CP-element group 382:  transition  input  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	374 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	412 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_update_completed_
      -- CP-element group 382: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_Update/$exit
      -- CP-element group 382: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_Update/ca
      -- 
    ca_2872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1225_inst_ack_1, ack => convTranspose_CP_34_elements(382)); -- 
    -- CP-element group 383:  transition  input  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	378 
    -- CP-element group 383: successors 
    -- CP-element group 383:  members (3) 
      -- CP-element group 383: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_sample_completed_
      -- CP-element group 383: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_Sample/$exit
      -- CP-element group 383: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_Sample/ra
      -- 
    ra_2881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1235_inst_ack_0, ack => convTranspose_CP_34_elements(383)); -- 
    -- CP-element group 384:  transition  input  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	374 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	409 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_update_completed_
      -- CP-element group 384: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_Update/$exit
      -- CP-element group 384: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_Update/ca
      -- 
    ca_2886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1235_inst_ack_1, ack => convTranspose_CP_34_elements(384)); -- 
    -- CP-element group 385:  transition  input  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	378 
    -- CP-element group 385: successors 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_sample_completed_
      -- CP-element group 385: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_Sample/$exit
      -- CP-element group 385: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_Sample/ra
      -- 
    ra_2895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1245_inst_ack_0, ack => convTranspose_CP_34_elements(385)); -- 
    -- CP-element group 386:  transition  input  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	374 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	406 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_update_completed_
      -- CP-element group 386: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_Update/$exit
      -- CP-element group 386: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_Update/ca
      -- 
    ca_2900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1245_inst_ack_1, ack => convTranspose_CP_34_elements(386)); -- 
    -- CP-element group 387:  transition  input  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	378 
    -- CP-element group 387: successors 
    -- CP-element group 387:  members (3) 
      -- CP-element group 387: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_sample_completed_
      -- CP-element group 387: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_Sample/$exit
      -- CP-element group 387: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_Sample/ra
      -- 
    ra_2909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1255_inst_ack_0, ack => convTranspose_CP_34_elements(387)); -- 
    -- CP-element group 388:  transition  input  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	374 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	403 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_update_completed_
      -- CP-element group 388: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_Update/$exit
      -- CP-element group 388: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_Update/ca
      -- 
    ca_2914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1255_inst_ack_1, ack => convTranspose_CP_34_elements(388)); -- 
    -- CP-element group 389:  transition  input  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	378 
    -- CP-element group 389: successors 
    -- CP-element group 389:  members (3) 
      -- CP-element group 389: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_sample_completed_
      -- CP-element group 389: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_Sample/$exit
      -- CP-element group 389: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_Sample/ra
      -- 
    ra_2923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1265_inst_ack_0, ack => convTranspose_CP_34_elements(389)); -- 
    -- CP-element group 390:  transition  input  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	374 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	400 
    -- CP-element group 390:  members (3) 
      -- CP-element group 390: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_update_completed_
      -- CP-element group 390: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_Update/$exit
      -- CP-element group 390: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_Update/ca
      -- 
    ca_2928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1265_inst_ack_1, ack => convTranspose_CP_34_elements(390)); -- 
    -- CP-element group 391:  transition  input  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	378 
    -- CP-element group 391: successors 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_sample_completed_
      -- CP-element group 391: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_Sample/$exit
      -- CP-element group 391: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_Sample/ra
      -- 
    ra_2937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1275_inst_ack_0, ack => convTranspose_CP_34_elements(391)); -- 
    -- CP-element group 392:  transition  input  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	374 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	397 
    -- CP-element group 392:  members (3) 
      -- CP-element group 392: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_update_completed_
      -- CP-element group 392: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_Update/$exit
      -- CP-element group 392: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_Update/ca
      -- 
    ca_2942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1275_inst_ack_1, ack => convTranspose_CP_34_elements(392)); -- 
    -- CP-element group 393:  transition  input  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	378 
    -- CP-element group 393: successors 
    -- CP-element group 393:  members (3) 
      -- CP-element group 393: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_sample_completed_
      -- CP-element group 393: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_Sample/$exit
      -- CP-element group 393: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_Sample/ra
      -- 
    ra_2951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1285_inst_ack_0, ack => convTranspose_CP_34_elements(393)); -- 
    -- CP-element group 394:  transition  input  output  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	374 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	395 
    -- CP-element group 394:  members (6) 
      -- CP-element group 394: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_update_completed_
      -- CP-element group 394: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_Update/$exit
      -- CP-element group 394: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_Update/ca
      -- CP-element group 394: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_sample_start_
      -- CP-element group 394: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_Sample/$entry
      -- CP-element group 394: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_Sample/req
      -- 
    ca_2956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1285_inst_ack_1, ack => convTranspose_CP_34_elements(394)); -- 
    req_2964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(394), ack => WPIPE_ConvTranspose_output_pipe_1287_inst_req_0); -- 
    -- CP-element group 395:  transition  input  output  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	394 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	396 
    -- CP-element group 395:  members (6) 
      -- CP-element group 395: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_Update/req
      -- CP-element group 395: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_Update/$entry
      -- CP-element group 395: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_sample_completed_
      -- CP-element group 395: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_update_start_
      -- CP-element group 395: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_Sample/$exit
      -- CP-element group 395: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_Sample/ack
      -- 
    ack_2965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1287_inst_ack_0, ack => convTranspose_CP_34_elements(395)); -- 
    req_2969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(395), ack => WPIPE_ConvTranspose_output_pipe_1287_inst_req_1); -- 
    -- CP-element group 396:  transition  input  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	395 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	397 
    -- CP-element group 396:  members (3) 
      -- CP-element group 396: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_Update/$exit
      -- CP-element group 396: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_Update/ack
      -- CP-element group 396: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_update_completed_
      -- 
    ack_2970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1287_inst_ack_1, ack => convTranspose_CP_34_elements(396)); -- 
    -- CP-element group 397:  join  transition  output  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	392 
    -- CP-element group 397: 	396 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	398 
    -- CP-element group 397:  members (3) 
      -- CP-element group 397: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_sample_start_
      -- CP-element group 397: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_Sample/req
      -- CP-element group 397: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_Sample/$entry
      -- 
    req_2978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(397), ack => WPIPE_ConvTranspose_output_pipe_1290_inst_req_0); -- 
    convTranspose_cp_element_group_397: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_397"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(392) & convTranspose_CP_34_elements(396);
      gj_convTranspose_cp_element_group_397 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(397), clk => clk, reset => reset); --
    end block;
    -- CP-element group 398:  transition  input  output  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	397 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	399 
    -- CP-element group 398:  members (6) 
      -- CP-element group 398: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_Sample/$exit
      -- CP-element group 398: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_Sample/ack
      -- CP-element group 398: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_update_start_
      -- CP-element group 398: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_Update/$entry
      -- CP-element group 398: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_sample_completed_
      -- CP-element group 398: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_Update/req
      -- 
    ack_2979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 398_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1290_inst_ack_0, ack => convTranspose_CP_34_elements(398)); -- 
    req_2983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(398), ack => WPIPE_ConvTranspose_output_pipe_1290_inst_req_1); -- 
    -- CP-element group 399:  transition  input  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	398 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	400 
    -- CP-element group 399:  members (3) 
      -- CP-element group 399: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_Update/$exit
      -- CP-element group 399: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_update_completed_
      -- CP-element group 399: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_Update/ack
      -- 
    ack_2984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1290_inst_ack_1, ack => convTranspose_CP_34_elements(399)); -- 
    -- CP-element group 400:  join  transition  output  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	390 
    -- CP-element group 400: 	399 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	401 
    -- CP-element group 400:  members (3) 
      -- CP-element group 400: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_Sample/req
      -- CP-element group 400: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_Sample/$entry
      -- CP-element group 400: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_sample_start_
      -- 
    req_2992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(400), ack => WPIPE_ConvTranspose_output_pipe_1293_inst_req_0); -- 
    convTranspose_cp_element_group_400: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_400"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(390) & convTranspose_CP_34_elements(399);
      gj_convTranspose_cp_element_group_400 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(400), clk => clk, reset => reset); --
    end block;
    -- CP-element group 401:  transition  input  output  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	400 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	402 
    -- CP-element group 401:  members (6) 
      -- CP-element group 401: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_Update/req
      -- CP-element group 401: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_Update/$entry
      -- CP-element group 401: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_Sample/ack
      -- CP-element group 401: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_Sample/$exit
      -- CP-element group 401: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_update_start_
      -- CP-element group 401: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_sample_completed_
      -- 
    ack_2993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1293_inst_ack_0, ack => convTranspose_CP_34_elements(401)); -- 
    req_2997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(401), ack => WPIPE_ConvTranspose_output_pipe_1293_inst_req_1); -- 
    -- CP-element group 402:  transition  input  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	401 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	403 
    -- CP-element group 402:  members (3) 
      -- CP-element group 402: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_Update/ack
      -- CP-element group 402: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_Update/$exit
      -- CP-element group 402: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_update_completed_
      -- 
    ack_2998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 402_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1293_inst_ack_1, ack => convTranspose_CP_34_elements(402)); -- 
    -- CP-element group 403:  join  transition  output  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	388 
    -- CP-element group 403: 	402 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	404 
    -- CP-element group 403:  members (3) 
      -- CP-element group 403: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_Sample/req
      -- CP-element group 403: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_Sample/$entry
      -- CP-element group 403: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_sample_start_
      -- 
    req_3006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(403), ack => WPIPE_ConvTranspose_output_pipe_1296_inst_req_0); -- 
    convTranspose_cp_element_group_403: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_403"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(388) & convTranspose_CP_34_elements(402);
      gj_convTranspose_cp_element_group_403 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(403), clk => clk, reset => reset); --
    end block;
    -- CP-element group 404:  transition  input  output  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	403 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	405 
    -- CP-element group 404:  members (6) 
      -- CP-element group 404: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_Update/req
      -- CP-element group 404: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_Sample/ack
      -- CP-element group 404: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_Sample/$exit
      -- CP-element group 404: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_update_start_
      -- CP-element group 404: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_sample_completed_
      -- 
    ack_3007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1296_inst_ack_0, ack => convTranspose_CP_34_elements(404)); -- 
    req_3011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(404), ack => WPIPE_ConvTranspose_output_pipe_1296_inst_req_1); -- 
    -- CP-element group 405:  transition  input  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	404 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	406 
    -- CP-element group 405:  members (3) 
      -- CP-element group 405: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_Update/ack
      -- CP-element group 405: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_Update/$exit
      -- CP-element group 405: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_update_completed_
      -- 
    ack_3012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 405_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1296_inst_ack_1, ack => convTranspose_CP_34_elements(405)); -- 
    -- CP-element group 406:  join  transition  output  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	386 
    -- CP-element group 406: 	405 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	407 
    -- CP-element group 406:  members (3) 
      -- CP-element group 406: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_Sample/req
      -- CP-element group 406: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_Sample/$entry
      -- CP-element group 406: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_sample_start_
      -- 
    req_3020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(406), ack => WPIPE_ConvTranspose_output_pipe_1299_inst_req_0); -- 
    convTranspose_cp_element_group_406: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_406"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(386) & convTranspose_CP_34_elements(405);
      gj_convTranspose_cp_element_group_406 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(406), clk => clk, reset => reset); --
    end block;
    -- CP-element group 407:  transition  input  output  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	406 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	408 
    -- CP-element group 407:  members (6) 
      -- CP-element group 407: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_Update/req
      -- CP-element group 407: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_Sample/$exit
      -- CP-element group 407: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_Update/$entry
      -- CP-element group 407: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_Sample/ack
      -- CP-element group 407: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_update_start_
      -- CP-element group 407: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_sample_completed_
      -- 
    ack_3021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1299_inst_ack_0, ack => convTranspose_CP_34_elements(407)); -- 
    req_3025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(407), ack => WPIPE_ConvTranspose_output_pipe_1299_inst_req_1); -- 
    -- CP-element group 408:  transition  input  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	407 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	409 
    -- CP-element group 408:  members (3) 
      -- CP-element group 408: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_Update/ack
      -- CP-element group 408: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_Update/$exit
      -- CP-element group 408: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_update_completed_
      -- 
    ack_3026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 408_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1299_inst_ack_1, ack => convTranspose_CP_34_elements(408)); -- 
    -- CP-element group 409:  join  transition  output  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	384 
    -- CP-element group 409: 	408 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	410 
    -- CP-element group 409:  members (3) 
      -- CP-element group 409: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_Sample/req
      -- CP-element group 409: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_sample_start_
      -- CP-element group 409: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_Sample/$entry
      -- 
    req_3034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(409), ack => WPIPE_ConvTranspose_output_pipe_1302_inst_req_0); -- 
    convTranspose_cp_element_group_409: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_409"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(384) & convTranspose_CP_34_elements(408);
      gj_convTranspose_cp_element_group_409 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(409), clk => clk, reset => reset); --
    end block;
    -- CP-element group 410:  transition  input  output  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	409 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	411 
    -- CP-element group 410:  members (6) 
      -- CP-element group 410: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_Update/req
      -- CP-element group 410: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_sample_completed_
      -- CP-element group 410: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_update_start_
      -- CP-element group 410: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_Sample/$exit
      -- CP-element group 410: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_Sample/ack
      -- 
    ack_3035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1302_inst_ack_0, ack => convTranspose_CP_34_elements(410)); -- 
    req_3039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(410), ack => WPIPE_ConvTranspose_output_pipe_1302_inst_req_1); -- 
    -- CP-element group 411:  transition  input  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	410 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	412 
    -- CP-element group 411:  members (3) 
      -- CP-element group 411: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_Update/$exit
      -- CP-element group 411: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_update_completed_
      -- CP-element group 411: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_Update/ack
      -- 
    ack_3040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 411_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1302_inst_ack_1, ack => convTranspose_CP_34_elements(411)); -- 
    -- CP-element group 412:  join  transition  output  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	382 
    -- CP-element group 412: 	411 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	413 
    -- CP-element group 412:  members (3) 
      -- CP-element group 412: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_Sample/$entry
      -- CP-element group 412: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_sample_start_
      -- CP-element group 412: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_Sample/req
      -- 
    req_3048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(412), ack => WPIPE_ConvTranspose_output_pipe_1305_inst_req_0); -- 
    convTranspose_cp_element_group_412: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_412"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(382) & convTranspose_CP_34_elements(411);
      gj_convTranspose_cp_element_group_412 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(412), clk => clk, reset => reset); --
    end block;
    -- CP-element group 413:  transition  input  output  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	412 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	414 
    -- CP-element group 413:  members (6) 
      -- CP-element group 413: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_update_start_
      -- CP-element group 413: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_sample_completed_
      -- CP-element group 413: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_Update/req
      -- CP-element group 413: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_Update/$entry
      -- CP-element group 413: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_Sample/ack
      -- CP-element group 413: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_Sample/$exit
      -- 
    ack_3049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1305_inst_ack_0, ack => convTranspose_CP_34_elements(413)); -- 
    req_3053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(413), ack => WPIPE_ConvTranspose_output_pipe_1305_inst_req_1); -- 
    -- CP-element group 414:  transition  input  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	413 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	415 
    -- CP-element group 414:  members (3) 
      -- CP-element group 414: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_update_completed_
      -- CP-element group 414: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_Update/ack
      -- CP-element group 414: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_Update/$exit
      -- 
    ack_3054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 414_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1305_inst_ack_1, ack => convTranspose_CP_34_elements(414)); -- 
    -- CP-element group 415:  join  transition  output  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	380 
    -- CP-element group 415: 	414 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	416 
    -- CP-element group 415:  members (3) 
      -- CP-element group 415: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_Sample/req
      -- CP-element group 415: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_Sample/$entry
      -- CP-element group 415: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_sample_start_
      -- 
    req_3062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(415), ack => WPIPE_ConvTranspose_output_pipe_1308_inst_req_0); -- 
    convTranspose_cp_element_group_415: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_415"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(380) & convTranspose_CP_34_elements(414);
      gj_convTranspose_cp_element_group_415 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(415), clk => clk, reset => reset); --
    end block;
    -- CP-element group 416:  transition  input  output  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	415 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	417 
    -- CP-element group 416:  members (6) 
      -- CP-element group 416: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_Update/req
      -- CP-element group 416: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_Update/$entry
      -- CP-element group 416: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_Sample/ack
      -- CP-element group 416: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_Sample/$exit
      -- CP-element group 416: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_update_start_
      -- CP-element group 416: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_sample_completed_
      -- 
    ack_3063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1308_inst_ack_0, ack => convTranspose_CP_34_elements(416)); -- 
    req_3067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(416), ack => WPIPE_ConvTranspose_output_pipe_1308_inst_req_1); -- 
    -- CP-element group 417:  branch  transition  place  input  output  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	416 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	418 
    -- CP-element group 417: 	419 
    -- CP-element group 417:  members (13) 
      -- CP-element group 417: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310__exit__
      -- CP-element group 417: 	 branch_block_stmt_38/if_stmt_1312__entry__
      -- CP-element group 417: 	 branch_block_stmt_38/if_stmt_1312_else_link/$entry
      -- CP-element group 417: 	 branch_block_stmt_38/if_stmt_1312_if_link/$entry
      -- CP-element group 417: 	 branch_block_stmt_38/if_stmt_1312_eval_test/branch_req
      -- CP-element group 417: 	 branch_block_stmt_38/if_stmt_1312_eval_test/$exit
      -- CP-element group 417: 	 branch_block_stmt_38/if_stmt_1312_eval_test/$entry
      -- CP-element group 417: 	 branch_block_stmt_38/if_stmt_1312_dead_link/$entry
      -- CP-element group 417: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_Update/ack
      -- CP-element group 417: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_Update/$exit
      -- CP-element group 417: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_update_completed_
      -- CP-element group 417: 	 branch_block_stmt_38/R_cmp264505_1313_place
      -- CP-element group 417: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/$exit
      -- 
    ack_3068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1308_inst_ack_1, ack => convTranspose_CP_34_elements(417)); -- 
    branch_req_3076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(417), ack => if_stmt_1312_branch_req_0); -- 
    -- CP-element group 418:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	417 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	420 
    -- CP-element group 418: 	421 
    -- CP-element group 418:  members (18) 
      -- CP-element group 418: 	 branch_block_stmt_38/merge_stmt_1318__exit__
      -- CP-element group 418: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353__entry__
      -- CP-element group 418: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_Update/cr
      -- CP-element group 418: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_Update/$entry
      -- CP-element group 418: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_Sample/rr
      -- CP-element group 418: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_update_start_
      -- CP-element group 418: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/$entry
      -- CP-element group 418: 	 branch_block_stmt_38/if_stmt_1312_if_link/if_choice_transition
      -- CP-element group 418: 	 branch_block_stmt_38/if_stmt_1312_if_link/$exit
      -- CP-element group 418: 	 branch_block_stmt_38/forx_xend273_bbx_xnph
      -- CP-element group 418: 	 branch_block_stmt_38/forx_xend273_bbx_xnph_PhiReq/$entry
      -- CP-element group 418: 	 branch_block_stmt_38/forx_xend273_bbx_xnph_PhiReq/$exit
      -- CP-element group 418: 	 branch_block_stmt_38/merge_stmt_1318_PhiReqMerge
      -- CP-element group 418: 	 branch_block_stmt_38/merge_stmt_1318_PhiAck/$entry
      -- CP-element group 418: 	 branch_block_stmt_38/merge_stmt_1318_PhiAck/$exit
      -- CP-element group 418: 	 branch_block_stmt_38/merge_stmt_1318_PhiAck/dummy
      -- 
    if_choice_transition_3081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 418_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1312_branch_ack_1, ack => convTranspose_CP_34_elements(418)); -- 
    cr_3103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(418), ack => type_cast_1339_inst_req_1); -- 
    rr_3098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(418), ack => type_cast_1339_inst_req_0); -- 
    -- CP-element group 419:  transition  place  input  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	417 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	497 
    -- CP-element group 419:  members (5) 
      -- CP-element group 419: 	 branch_block_stmt_38/forx_xend273_forx_xend500
      -- CP-element group 419: 	 branch_block_stmt_38/if_stmt_1312_else_link/else_choice_transition
      -- CP-element group 419: 	 branch_block_stmt_38/if_stmt_1312_else_link/$exit
      -- CP-element group 419: 	 branch_block_stmt_38/forx_xend273_forx_xend500_PhiReq/$entry
      -- CP-element group 419: 	 branch_block_stmt_38/forx_xend273_forx_xend500_PhiReq/$exit
      -- 
    else_choice_transition_3085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1312_branch_ack_0, ack => convTranspose_CP_34_elements(419)); -- 
    -- CP-element group 420:  transition  input  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	418 
    -- CP-element group 420: successors 
    -- CP-element group 420:  members (3) 
      -- CP-element group 420: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_Sample/ra
      -- CP-element group 420: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_Sample/$exit
      -- CP-element group 420: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_sample_completed_
      -- 
    ra_3099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1339_inst_ack_0, ack => convTranspose_CP_34_elements(420)); -- 
    -- CP-element group 421:  transition  place  input  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	418 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	491 
    -- CP-element group 421:  members (9) 
      -- CP-element group 421: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353__exit__
      -- CP-element group 421: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427
      -- CP-element group 421: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_Update/ca
      -- CP-element group 421: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_Update/$exit
      -- CP-element group 421: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_update_completed_
      -- CP-element group 421: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/$exit
      -- CP-element group 421: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/$entry
      -- CP-element group 421: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1356/$entry
      -- CP-element group 421: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/$entry
      -- 
    ca_3104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1339_inst_ack_1, ack => convTranspose_CP_34_elements(421)); -- 
    -- CP-element group 422:  transition  input  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	496 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	467 
    -- CP-element group 422:  members (3) 
      -- CP-element group 422: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_final_index_sum_regn_sample_complete
      -- CP-element group 422: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_final_index_sum_regn_Sample/ack
      -- CP-element group 422: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_final_index_sum_regn_Sample/$exit
      -- 
    ack_3133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 422_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1368_index_offset_ack_0, ack => convTranspose_CP_34_elements(422)); -- 
    -- CP-element group 423:  transition  input  output  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	496 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	424 
    -- CP-element group 423:  members (11) 
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_sample_start_
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_root_address_calculated
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_offset_calculated
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_request/req
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_request/$entry
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_base_plus_offset/sum_rename_ack
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_base_plus_offset/sum_rename_req
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_base_plus_offset/$exit
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_base_plus_offset/$entry
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_final_index_sum_regn_Update/ack
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_final_index_sum_regn_Update/$exit
      -- 
    ack_3138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 423_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1368_index_offset_ack_1, ack => convTranspose_CP_34_elements(423)); -- 
    req_3147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(423), ack => addr_of_1369_final_reg_req_0); -- 
    -- CP-element group 424:  transition  input  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	423 
    -- CP-element group 424: successors 
    -- CP-element group 424:  members (3) 
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_sample_completed_
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_request/ack
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_request/$exit
      -- 
    ack_3148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1369_final_reg_ack_0, ack => convTranspose_CP_34_elements(424)); -- 
    -- CP-element group 425:  join  fork  transition  input  output  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	496 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	426 
    -- CP-element group 425:  members (24) 
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_update_completed_
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Sample/word_access_start/word_0/rr
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Sample/word_access_start/word_0/$entry
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Sample/word_access_start/$entry
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Sample/$entry
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_word_addrgen/root_register_ack
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_word_addrgen/root_register_req
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_word_addrgen/$exit
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_word_addrgen/$entry
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_base_plus_offset/sum_rename_ack
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_base_plus_offset/sum_rename_req
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_base_plus_offset/$exit
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_base_plus_offset/$entry
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_base_addr_resize/base_resize_ack
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_base_addr_resize/base_resize_req
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_base_addr_resize/$exit
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_base_addr_resize/$entry
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_base_address_resized
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_root_address_calculated
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_word_address_calculated
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_base_address_calculated
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_sample_start_
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_complete/ack
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_complete/$exit
      -- 
    ack_3153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1369_final_reg_ack_1, ack => convTranspose_CP_34_elements(425)); -- 
    rr_3186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(425), ack => ptr_deref_1373_load_0_req_0); -- 
    -- CP-element group 426:  transition  input  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	425 
    -- CP-element group 426: successors 
    -- CP-element group 426:  members (5) 
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Sample/word_access_start/word_0/ra
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Sample/word_access_start/word_0/$exit
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Sample/word_access_start/$exit
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Sample/$exit
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_sample_completed_
      -- 
    ra_3187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 426_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1373_load_0_ack_0, ack => convTranspose_CP_34_elements(426)); -- 
    -- CP-element group 427:  fork  transition  input  output  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	496 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	428 
    -- CP-element group 427: 	430 
    -- CP-element group 427: 	432 
    -- CP-element group 427: 	434 
    -- CP-element group 427: 	436 
    -- CP-element group 427: 	438 
    -- CP-element group 427: 	440 
    -- CP-element group 427: 	442 
    -- CP-element group 427:  members (33) 
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/word_access_complete/word_0/$exit
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/ptr_deref_1373_Merge/$entry
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/word_access_complete/word_0/ca
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_Sample/rr
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/word_access_complete/$exit
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/$exit
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_Sample/rr
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_Sample/rr
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_Sample/rr
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_Sample/rr
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_update_completed_
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_Sample/rr
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_Sample/rr
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/ptr_deref_1373_Merge/merge_ack
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/ptr_deref_1373_Merge/merge_req
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/ptr_deref_1373_Merge/$exit
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_Sample/rr
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_sample_start_
      -- 
    ca_3198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 427_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1373_load_0_ack_1, ack => convTranspose_CP_34_elements(427)); -- 
    rr_3211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(427), ack => type_cast_1377_inst_req_0); -- 
    rr_3225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(427), ack => type_cast_1387_inst_req_0); -- 
    rr_3239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(427), ack => type_cast_1397_inst_req_0); -- 
    rr_3253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(427), ack => type_cast_1407_inst_req_0); -- 
    rr_3267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(427), ack => type_cast_1417_inst_req_0); -- 
    rr_3281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(427), ack => type_cast_1427_inst_req_0); -- 
    rr_3295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(427), ack => type_cast_1437_inst_req_0); -- 
    rr_3309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(427), ack => type_cast_1447_inst_req_0); -- 
    -- CP-element group 428:  transition  input  bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	427 
    -- CP-element group 428: successors 
    -- CP-element group 428:  members (3) 
      -- CP-element group 428: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_Sample/ra
      -- CP-element group 428: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_Sample/$exit
      -- CP-element group 428: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_sample_completed_
      -- 
    ra_3212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1377_inst_ack_0, ack => convTranspose_CP_34_elements(428)); -- 
    -- CP-element group 429:  transition  input  bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	496 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	464 
    -- CP-element group 429:  members (3) 
      -- CP-element group 429: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_Update/ca
      -- CP-element group 429: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_Update/$exit
      -- CP-element group 429: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_update_completed_
      -- 
    ca_3217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1377_inst_ack_1, ack => convTranspose_CP_34_elements(429)); -- 
    -- CP-element group 430:  transition  input  bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	427 
    -- CP-element group 430: successors 
    -- CP-element group 430:  members (3) 
      -- CP-element group 430: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_Sample/ra
      -- CP-element group 430: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_Sample/$exit
      -- CP-element group 430: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_sample_completed_
      -- 
    ra_3226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 430_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1387_inst_ack_0, ack => convTranspose_CP_34_elements(430)); -- 
    -- CP-element group 431:  transition  input  bypass 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	496 
    -- CP-element group 431: successors 
    -- CP-element group 431: 	461 
    -- CP-element group 431:  members (3) 
      -- CP-element group 431: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_Update/ca
      -- CP-element group 431: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_Update/$exit
      -- CP-element group 431: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_update_completed_
      -- 
    ca_3231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 431_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1387_inst_ack_1, ack => convTranspose_CP_34_elements(431)); -- 
    -- CP-element group 432:  transition  input  bypass 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	427 
    -- CP-element group 432: successors 
    -- CP-element group 432:  members (3) 
      -- CP-element group 432: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_sample_completed_
      -- CP-element group 432: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_Sample/$exit
      -- CP-element group 432: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_Sample/ra
      -- 
    ra_3240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1397_inst_ack_0, ack => convTranspose_CP_34_elements(432)); -- 
    -- CP-element group 433:  transition  input  bypass 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	496 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	458 
    -- CP-element group 433:  members (3) 
      -- CP-element group 433: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_update_completed_
      -- CP-element group 433: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_Update/ca
      -- CP-element group 433: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_Update/$exit
      -- 
    ca_3245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1397_inst_ack_1, ack => convTranspose_CP_34_elements(433)); -- 
    -- CP-element group 434:  transition  input  bypass 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	427 
    -- CP-element group 434: successors 
    -- CP-element group 434:  members (3) 
      -- CP-element group 434: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_Sample/ra
      -- CP-element group 434: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_Sample/$exit
      -- CP-element group 434: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_sample_completed_
      -- 
    ra_3254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 434_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1407_inst_ack_0, ack => convTranspose_CP_34_elements(434)); -- 
    -- CP-element group 435:  transition  input  bypass 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	496 
    -- CP-element group 435: successors 
    -- CP-element group 435: 	455 
    -- CP-element group 435:  members (3) 
      -- CP-element group 435: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_Update/ca
      -- CP-element group 435: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_Update/$exit
      -- CP-element group 435: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_update_completed_
      -- 
    ca_3259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1407_inst_ack_1, ack => convTranspose_CP_34_elements(435)); -- 
    -- CP-element group 436:  transition  input  bypass 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	427 
    -- CP-element group 436: successors 
    -- CP-element group 436:  members (3) 
      -- CP-element group 436: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_Sample/$exit
      -- CP-element group 436: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_Sample/ra
      -- CP-element group 436: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_sample_completed_
      -- 
    ra_3268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1417_inst_ack_0, ack => convTranspose_CP_34_elements(436)); -- 
    -- CP-element group 437:  transition  input  bypass 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	496 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	452 
    -- CP-element group 437:  members (3) 
      -- CP-element group 437: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_Update/ca
      -- CP-element group 437: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_update_completed_
      -- CP-element group 437: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_Update/$exit
      -- 
    ca_3273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 437_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1417_inst_ack_1, ack => convTranspose_CP_34_elements(437)); -- 
    -- CP-element group 438:  transition  input  bypass 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	427 
    -- CP-element group 438: successors 
    -- CP-element group 438:  members (3) 
      -- CP-element group 438: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_Sample/ra
      -- CP-element group 438: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_Sample/$exit
      -- CP-element group 438: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_sample_completed_
      -- 
    ra_3282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 438_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1427_inst_ack_0, ack => convTranspose_CP_34_elements(438)); -- 
    -- CP-element group 439:  transition  input  bypass 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	496 
    -- CP-element group 439: successors 
    -- CP-element group 439: 	449 
    -- CP-element group 439:  members (3) 
      -- CP-element group 439: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_Update/ca
      -- CP-element group 439: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_Update/$exit
      -- CP-element group 439: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_update_completed_
      -- 
    ca_3287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 439_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1427_inst_ack_1, ack => convTranspose_CP_34_elements(439)); -- 
    -- CP-element group 440:  transition  input  bypass 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	427 
    -- CP-element group 440: successors 
    -- CP-element group 440:  members (3) 
      -- CP-element group 440: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_sample_completed_
      -- CP-element group 440: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_Sample/ra
      -- CP-element group 440: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_Sample/$exit
      -- 
    ra_3296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 440_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1437_inst_ack_0, ack => convTranspose_CP_34_elements(440)); -- 
    -- CP-element group 441:  transition  input  bypass 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	496 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	446 
    -- CP-element group 441:  members (3) 
      -- CP-element group 441: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_Update/ca
      -- CP-element group 441: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_Update/$exit
      -- CP-element group 441: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_update_completed_
      -- 
    ca_3301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 441_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1437_inst_ack_1, ack => convTranspose_CP_34_elements(441)); -- 
    -- CP-element group 442:  transition  input  bypass 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	427 
    -- CP-element group 442: successors 
    -- CP-element group 442:  members (3) 
      -- CP-element group 442: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_Sample/ra
      -- CP-element group 442: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_Sample/$exit
      -- CP-element group 442: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_sample_completed_
      -- 
    ra_3310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 442_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1447_inst_ack_0, ack => convTranspose_CP_34_elements(442)); -- 
    -- CP-element group 443:  transition  input  output  bypass 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	496 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	444 
    -- CP-element group 443:  members (6) 
      -- CP-element group 443: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_Sample/req
      -- CP-element group 443: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_Sample/$entry
      -- CP-element group 443: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_sample_start_
      -- CP-element group 443: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_Update/ca
      -- CP-element group 443: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_Update/$exit
      -- CP-element group 443: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_update_completed_
      -- 
    ca_3315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 443_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1447_inst_ack_1, ack => convTranspose_CP_34_elements(443)); -- 
    req_3323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(443), ack => WPIPE_ConvTranspose_output_pipe_1449_inst_req_0); -- 
    -- CP-element group 444:  transition  input  output  bypass 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	443 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	445 
    -- CP-element group 444:  members (6) 
      -- CP-element group 444: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_Update/req
      -- CP-element group 444: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_Update/$entry
      -- CP-element group 444: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_Sample/ack
      -- CP-element group 444: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_Sample/$exit
      -- CP-element group 444: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_update_start_
      -- CP-element group 444: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_sample_completed_
      -- 
    ack_3324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1449_inst_ack_0, ack => convTranspose_CP_34_elements(444)); -- 
    req_3328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(444), ack => WPIPE_ConvTranspose_output_pipe_1449_inst_req_1); -- 
    -- CP-element group 445:  transition  input  bypass 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	444 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	446 
    -- CP-element group 445:  members (3) 
      -- CP-element group 445: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_Update/ack
      -- CP-element group 445: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_Update/$exit
      -- CP-element group 445: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_update_completed_
      -- 
    ack_3329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 445_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1449_inst_ack_1, ack => convTranspose_CP_34_elements(445)); -- 
    -- CP-element group 446:  join  transition  output  bypass 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	441 
    -- CP-element group 446: 	445 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	447 
    -- CP-element group 446:  members (3) 
      -- CP-element group 446: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_Sample/req
      -- CP-element group 446: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_Sample/$entry
      -- CP-element group 446: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_sample_start_
      -- 
    req_3337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(446), ack => WPIPE_ConvTranspose_output_pipe_1452_inst_req_0); -- 
    convTranspose_cp_element_group_446: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_446"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(441) & convTranspose_CP_34_elements(445);
      gj_convTranspose_cp_element_group_446 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(446), clk => clk, reset => reset); --
    end block;
    -- CP-element group 447:  transition  input  output  bypass 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	446 
    -- CP-element group 447: successors 
    -- CP-element group 447: 	448 
    -- CP-element group 447:  members (6) 
      -- CP-element group 447: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_Update/req
      -- CP-element group 447: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_Update/$entry
      -- CP-element group 447: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_Sample/ack
      -- CP-element group 447: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_Sample/$exit
      -- CP-element group 447: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_update_start_
      -- CP-element group 447: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_sample_completed_
      -- 
    ack_3338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1452_inst_ack_0, ack => convTranspose_CP_34_elements(447)); -- 
    req_3342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(447), ack => WPIPE_ConvTranspose_output_pipe_1452_inst_req_1); -- 
    -- CP-element group 448:  transition  input  bypass 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	447 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	449 
    -- CP-element group 448:  members (3) 
      -- CP-element group 448: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_Update/ack
      -- CP-element group 448: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_Update/$exit
      -- CP-element group 448: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_update_completed_
      -- 
    ack_3343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 448_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1452_inst_ack_1, ack => convTranspose_CP_34_elements(448)); -- 
    -- CP-element group 449:  join  transition  output  bypass 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	439 
    -- CP-element group 449: 	448 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	450 
    -- CP-element group 449:  members (3) 
      -- CP-element group 449: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_sample_start_
      -- CP-element group 449: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_Sample/req
      -- CP-element group 449: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_Sample/$entry
      -- 
    req_3351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(449), ack => WPIPE_ConvTranspose_output_pipe_1455_inst_req_0); -- 
    convTranspose_cp_element_group_449: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_449"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(439) & convTranspose_CP_34_elements(448);
      gj_convTranspose_cp_element_group_449 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(449), clk => clk, reset => reset); --
    end block;
    -- CP-element group 450:  transition  input  output  bypass 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	449 
    -- CP-element group 450: successors 
    -- CP-element group 450: 	451 
    -- CP-element group 450:  members (6) 
      -- CP-element group 450: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_update_start_
      -- CP-element group 450: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_Update/req
      -- CP-element group 450: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_sample_completed_
      -- CP-element group 450: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_Update/$entry
      -- CP-element group 450: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_Sample/ack
      -- CP-element group 450: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_Sample/$exit
      -- 
    ack_3352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 450_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1455_inst_ack_0, ack => convTranspose_CP_34_elements(450)); -- 
    req_3356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(450), ack => WPIPE_ConvTranspose_output_pipe_1455_inst_req_1); -- 
    -- CP-element group 451:  transition  input  bypass 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	450 
    -- CP-element group 451: successors 
    -- CP-element group 451: 	452 
    -- CP-element group 451:  members (3) 
      -- CP-element group 451: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_Update/ack
      -- CP-element group 451: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_Update/$exit
      -- CP-element group 451: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_update_completed_
      -- 
    ack_3357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 451_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1455_inst_ack_1, ack => convTranspose_CP_34_elements(451)); -- 
    -- CP-element group 452:  join  transition  output  bypass 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	437 
    -- CP-element group 452: 	451 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	453 
    -- CP-element group 452:  members (3) 
      -- CP-element group 452: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_Sample/req
      -- CP-element group 452: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_sample_start_
      -- 
    req_3365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(452), ack => WPIPE_ConvTranspose_output_pipe_1458_inst_req_0); -- 
    convTranspose_cp_element_group_452: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_452"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(437) & convTranspose_CP_34_elements(451);
      gj_convTranspose_cp_element_group_452 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(452), clk => clk, reset => reset); --
    end block;
    -- CP-element group 453:  transition  input  output  bypass 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	452 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	454 
    -- CP-element group 453:  members (6) 
      -- CP-element group 453: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_Update/req
      -- CP-element group 453: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_Update/$entry
      -- CP-element group 453: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_Sample/ack
      -- CP-element group 453: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_Sample/$exit
      -- CP-element group 453: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_update_start_
      -- CP-element group 453: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_sample_completed_
      -- 
    ack_3366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 453_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1458_inst_ack_0, ack => convTranspose_CP_34_elements(453)); -- 
    req_3370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(453), ack => WPIPE_ConvTranspose_output_pipe_1458_inst_req_1); -- 
    -- CP-element group 454:  transition  input  bypass 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	453 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	455 
    -- CP-element group 454:  members (3) 
      -- CP-element group 454: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_Update/ack
      -- CP-element group 454: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_Update/$exit
      -- CP-element group 454: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_update_completed_
      -- 
    ack_3371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 454_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1458_inst_ack_1, ack => convTranspose_CP_34_elements(454)); -- 
    -- CP-element group 455:  join  transition  output  bypass 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	435 
    -- CP-element group 455: 	454 
    -- CP-element group 455: successors 
    -- CP-element group 455: 	456 
    -- CP-element group 455:  members (3) 
      -- CP-element group 455: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_Sample/$entry
      -- CP-element group 455: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_sample_start_
      -- CP-element group 455: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_Sample/req
      -- 
    req_3379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(455), ack => WPIPE_ConvTranspose_output_pipe_1461_inst_req_0); -- 
    convTranspose_cp_element_group_455: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_455"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(435) & convTranspose_CP_34_elements(454);
      gj_convTranspose_cp_element_group_455 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(455), clk => clk, reset => reset); --
    end block;
    -- CP-element group 456:  transition  input  output  bypass 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	455 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	457 
    -- CP-element group 456:  members (6) 
      -- CP-element group 456: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_update_start_
      -- CP-element group 456: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_sample_completed_
      -- CP-element group 456: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_Sample/$exit
      -- CP-element group 456: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_Sample/ack
      -- CP-element group 456: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_Update/$entry
      -- CP-element group 456: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_Update/req
      -- 
    ack_3380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 456_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1461_inst_ack_0, ack => convTranspose_CP_34_elements(456)); -- 
    req_3384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(456), ack => WPIPE_ConvTranspose_output_pipe_1461_inst_req_1); -- 
    -- CP-element group 457:  transition  input  bypass 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	456 
    -- CP-element group 457: successors 
    -- CP-element group 457: 	458 
    -- CP-element group 457:  members (3) 
      -- CP-element group 457: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_update_completed_
      -- CP-element group 457: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_Update/$exit
      -- CP-element group 457: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_Update/ack
      -- 
    ack_3385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 457_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1461_inst_ack_1, ack => convTranspose_CP_34_elements(457)); -- 
    -- CP-element group 458:  join  transition  output  bypass 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	433 
    -- CP-element group 458: 	457 
    -- CP-element group 458: successors 
    -- CP-element group 458: 	459 
    -- CP-element group 458:  members (3) 
      -- CP-element group 458: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_sample_start_
      -- CP-element group 458: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_Sample/$entry
      -- CP-element group 458: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_Sample/req
      -- 
    req_3393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(458), ack => WPIPE_ConvTranspose_output_pipe_1464_inst_req_0); -- 
    convTranspose_cp_element_group_458: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_458"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(433) & convTranspose_CP_34_elements(457);
      gj_convTranspose_cp_element_group_458 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(458), clk => clk, reset => reset); --
    end block;
    -- CP-element group 459:  transition  input  output  bypass 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	458 
    -- CP-element group 459: successors 
    -- CP-element group 459: 	460 
    -- CP-element group 459:  members (6) 
      -- CP-element group 459: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_sample_completed_
      -- CP-element group 459: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_update_start_
      -- CP-element group 459: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_Sample/$exit
      -- CP-element group 459: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_Sample/ack
      -- CP-element group 459: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_Update/$entry
      -- CP-element group 459: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_Update/req
      -- 
    ack_3394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 459_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1464_inst_ack_0, ack => convTranspose_CP_34_elements(459)); -- 
    req_3398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(459), ack => WPIPE_ConvTranspose_output_pipe_1464_inst_req_1); -- 
    -- CP-element group 460:  transition  input  bypass 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	459 
    -- CP-element group 460: successors 
    -- CP-element group 460: 	461 
    -- CP-element group 460:  members (3) 
      -- CP-element group 460: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_update_completed_
      -- CP-element group 460: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_Update/$exit
      -- CP-element group 460: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_Update/ack
      -- 
    ack_3399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 460_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1464_inst_ack_1, ack => convTranspose_CP_34_elements(460)); -- 
    -- CP-element group 461:  join  transition  output  bypass 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	431 
    -- CP-element group 461: 	460 
    -- CP-element group 461: successors 
    -- CP-element group 461: 	462 
    -- CP-element group 461:  members (3) 
      -- CP-element group 461: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_sample_start_
      -- CP-element group 461: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_Sample/$entry
      -- CP-element group 461: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_Sample/req
      -- 
    req_3407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(461), ack => WPIPE_ConvTranspose_output_pipe_1467_inst_req_0); -- 
    convTranspose_cp_element_group_461: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_461"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(431) & convTranspose_CP_34_elements(460);
      gj_convTranspose_cp_element_group_461 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(461), clk => clk, reset => reset); --
    end block;
    -- CP-element group 462:  transition  input  output  bypass 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	461 
    -- CP-element group 462: successors 
    -- CP-element group 462: 	463 
    -- CP-element group 462:  members (6) 
      -- CP-element group 462: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_sample_completed_
      -- CP-element group 462: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_update_start_
      -- CP-element group 462: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_Sample/$exit
      -- CP-element group 462: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_Sample/ack
      -- CP-element group 462: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_Update/$entry
      -- CP-element group 462: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_Update/req
      -- 
    ack_3408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 462_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1467_inst_ack_0, ack => convTranspose_CP_34_elements(462)); -- 
    req_3412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(462), ack => WPIPE_ConvTranspose_output_pipe_1467_inst_req_1); -- 
    -- CP-element group 463:  transition  input  bypass 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	462 
    -- CP-element group 463: successors 
    -- CP-element group 463: 	464 
    -- CP-element group 463:  members (3) 
      -- CP-element group 463: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_update_completed_
      -- CP-element group 463: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_Update/$exit
      -- CP-element group 463: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_Update/ack
      -- 
    ack_3413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 463_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1467_inst_ack_1, ack => convTranspose_CP_34_elements(463)); -- 
    -- CP-element group 464:  join  transition  output  bypass 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	429 
    -- CP-element group 464: 	463 
    -- CP-element group 464: successors 
    -- CP-element group 464: 	465 
    -- CP-element group 464:  members (3) 
      -- CP-element group 464: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_sample_start_
      -- CP-element group 464: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_Sample/$entry
      -- CP-element group 464: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_Sample/req
      -- 
    req_3421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(464), ack => WPIPE_ConvTranspose_output_pipe_1470_inst_req_0); -- 
    convTranspose_cp_element_group_464: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_464"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(429) & convTranspose_CP_34_elements(463);
      gj_convTranspose_cp_element_group_464 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(464), clk => clk, reset => reset); --
    end block;
    -- CP-element group 465:  transition  input  output  bypass 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	464 
    -- CP-element group 465: successors 
    -- CP-element group 465: 	466 
    -- CP-element group 465:  members (6) 
      -- CP-element group 465: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_sample_completed_
      -- CP-element group 465: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_update_start_
      -- CP-element group 465: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_Sample/$exit
      -- CP-element group 465: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_Sample/ack
      -- CP-element group 465: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_Update/$entry
      -- CP-element group 465: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_Update/req
      -- 
    ack_3422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 465_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1470_inst_ack_0, ack => convTranspose_CP_34_elements(465)); -- 
    req_3426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(465), ack => WPIPE_ConvTranspose_output_pipe_1470_inst_req_1); -- 
    -- CP-element group 466:  transition  input  bypass 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	465 
    -- CP-element group 466: successors 
    -- CP-element group 466: 	467 
    -- CP-element group 466:  members (3) 
      -- CP-element group 466: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_update_completed_
      -- CP-element group 466: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_Update/$exit
      -- CP-element group 466: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_Update/ack
      -- 
    ack_3427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 466_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1470_inst_ack_1, ack => convTranspose_CP_34_elements(466)); -- 
    -- CP-element group 467:  branch  join  transition  place  output  bypass 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	422 
    -- CP-element group 467: 	466 
    -- CP-element group 467: successors 
    -- CP-element group 467: 	468 
    -- CP-element group 467: 	469 
    -- CP-element group 467:  members (10) 
      -- CP-element group 467: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483__exit__
      -- CP-element group 467: 	 branch_block_stmt_38/if_stmt_1484__entry__
      -- CP-element group 467: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/$exit
      -- CP-element group 467: 	 branch_block_stmt_38/if_stmt_1484_dead_link/$entry
      -- CP-element group 467: 	 branch_block_stmt_38/if_stmt_1484_eval_test/$entry
      -- CP-element group 467: 	 branch_block_stmt_38/if_stmt_1484_eval_test/$exit
      -- CP-element group 467: 	 branch_block_stmt_38/if_stmt_1484_eval_test/branch_req
      -- CP-element group 467: 	 branch_block_stmt_38/R_exitcond1_1485_place
      -- CP-element group 467: 	 branch_block_stmt_38/if_stmt_1484_if_link/$entry
      -- CP-element group 467: 	 branch_block_stmt_38/if_stmt_1484_else_link/$entry
      -- 
    branch_req_3435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(467), ack => if_stmt_1484_branch_req_0); -- 
    convTranspose_cp_element_group_467: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_467"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(422) & convTranspose_CP_34_elements(466);
      gj_convTranspose_cp_element_group_467 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(467), clk => clk, reset => reset); --
    end block;
    -- CP-element group 468:  merge  transition  place  input  bypass 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: 	467 
    -- CP-element group 468: successors 
    -- CP-element group 468: 	497 
    -- CP-element group 468:  members (13) 
      -- CP-element group 468: 	 branch_block_stmt_38/merge_stmt_1490__exit__
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xend500x_xloopexit_forx_xend500
      -- CP-element group 468: 	 branch_block_stmt_38/if_stmt_1484_if_link/$exit
      -- CP-element group 468: 	 branch_block_stmt_38/if_stmt_1484_if_link/if_choice_transition
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xbody427_forx_xend500x_xloopexit
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xbody427_forx_xend500x_xloopexit_PhiReq/$entry
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xbody427_forx_xend500x_xloopexit_PhiReq/$exit
      -- CP-element group 468: 	 branch_block_stmt_38/merge_stmt_1490_PhiReqMerge
      -- CP-element group 468: 	 branch_block_stmt_38/merge_stmt_1490_PhiAck/$entry
      -- CP-element group 468: 	 branch_block_stmt_38/merge_stmt_1490_PhiAck/$exit
      -- CP-element group 468: 	 branch_block_stmt_38/merge_stmt_1490_PhiAck/dummy
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xend500x_xloopexit_forx_xend500_PhiReq/$entry
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xend500x_xloopexit_forx_xend500_PhiReq/$exit
      -- 
    if_choice_transition_3440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 468_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1484_branch_ack_1, ack => convTranspose_CP_34_elements(468)); -- 
    -- CP-element group 469:  fork  transition  place  input  output  bypass 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	467 
    -- CP-element group 469: successors 
    -- CP-element group 469: 	492 
    -- CP-element group 469: 	493 
    -- CP-element group 469:  members (12) 
      -- CP-element group 469: 	 branch_block_stmt_38/if_stmt_1484_else_link/$exit
      -- CP-element group 469: 	 branch_block_stmt_38/if_stmt_1484_else_link/else_choice_transition
      -- CP-element group 469: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427
      -- CP-element group 469: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/$entry
      -- CP-element group 469: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/$entry
      -- CP-element group 469: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/$entry
      -- CP-element group 469: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/$entry
      -- CP-element group 469: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/SplitProtocol/$entry
      -- CP-element group 469: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/SplitProtocol/Sample/$entry
      -- CP-element group 469: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/SplitProtocol/Sample/rr
      -- CP-element group 469: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/SplitProtocol/Update/$entry
      -- CP-element group 469: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 469_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1484_branch_ack_0, ack => convTranspose_CP_34_elements(469)); -- 
    rr_3719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(469), ack => type_cast_1362_inst_req_0); -- 
    cr_3724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(469), ack => type_cast_1362_inst_req_1); -- 
    -- CP-element group 470:  merge  branch  transition  place  output  bypass 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	165 
    -- CP-element group 470: 	120 
    -- CP-element group 470: successors 
    -- CP-element group 470: 	121 
    -- CP-element group 470: 	122 
    -- CP-element group 470:  members (17) 
      -- CP-element group 470: 	 branch_block_stmt_38/merge_stmt_429__exit__
      -- CP-element group 470: 	 branch_block_stmt_38/assign_stmt_435__entry__
      -- CP-element group 470: 	 branch_block_stmt_38/assign_stmt_435__exit__
      -- CP-element group 470: 	 branch_block_stmt_38/if_stmt_436__entry__
      -- CP-element group 470: 	 branch_block_stmt_38/assign_stmt_435/$entry
      -- CP-element group 470: 	 branch_block_stmt_38/assign_stmt_435/$exit
      -- CP-element group 470: 	 branch_block_stmt_38/if_stmt_436_dead_link/$entry
      -- CP-element group 470: 	 branch_block_stmt_38/if_stmt_436_eval_test/$entry
      -- CP-element group 470: 	 branch_block_stmt_38/if_stmt_436_eval_test/$exit
      -- CP-element group 470: 	 branch_block_stmt_38/if_stmt_436_eval_test/branch_req
      -- CP-element group 470: 	 branch_block_stmt_38/R_cmp194509_437_place
      -- CP-element group 470: 	 branch_block_stmt_38/if_stmt_436_if_link/$entry
      -- CP-element group 470: 	 branch_block_stmt_38/if_stmt_436_else_link/$entry
      -- CP-element group 470: 	 branch_block_stmt_38/merge_stmt_429_PhiReqMerge
      -- CP-element group 470: 	 branch_block_stmt_38/merge_stmt_429_PhiAck/$entry
      -- CP-element group 470: 	 branch_block_stmt_38/merge_stmt_429_PhiAck/$exit
      -- CP-element group 470: 	 branch_block_stmt_38/merge_stmt_429_PhiAck/dummy
      -- 
    branch_req_924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(470), ack => if_stmt_436_branch_req_0); -- 
    convTranspose_CP_34_elements(470) <= OrReduce(convTranspose_CP_34_elements(165) & convTranspose_CP_34_elements(120));
    -- CP-element group 471:  transition  output  delay-element  bypass 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	124 
    -- CP-element group 471: successors 
    -- CP-element group 471: 	475 
    -- CP-element group 471:  members (5) 
      -- CP-element group 471: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/$exit
      -- CP-element group 471: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_474/$exit
      -- CP-element group 471: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/$exit
      -- CP-element group 471: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_478_konst_delay_trans
      -- CP-element group 471: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_req
      -- 
    phi_stmt_474_req_3492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_474_req_3492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(471), ack => phi_stmt_474_req_0); -- 
    -- Element group convTranspose_CP_34_elements(471) is a control-delay.
    cp_element_471_delay: control_delay_element  generic map(name => " 471_delay", delay_value => 1)  port map(req => convTranspose_CP_34_elements(124), ack => convTranspose_CP_34_elements(471), clk => clk, reset =>reset);
    -- CP-element group 472:  transition  input  bypass 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: 	166 
    -- CP-element group 472: successors 
    -- CP-element group 472: 	474 
    -- CP-element group 472:  members (2) 
      -- CP-element group 472: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Sample/$exit
      -- CP-element group 472: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Sample/ra
      -- 
    ra_3512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 472_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_480_inst_ack_0, ack => convTranspose_CP_34_elements(472)); -- 
    -- CP-element group 473:  transition  input  bypass 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	166 
    -- CP-element group 473: successors 
    -- CP-element group 473: 	474 
    -- CP-element group 473:  members (2) 
      -- CP-element group 473: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Update/$exit
      -- CP-element group 473: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Update/ca
      -- 
    ca_3517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 473_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_480_inst_ack_1, ack => convTranspose_CP_34_elements(473)); -- 
    -- CP-element group 474:  join  transition  output  bypass 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	472 
    -- CP-element group 474: 	473 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	475 
    -- CP-element group 474:  members (6) 
      -- CP-element group 474: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 474: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/$exit
      -- CP-element group 474: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/$exit
      -- CP-element group 474: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/$exit
      -- CP-element group 474: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/$exit
      -- CP-element group 474: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_req
      -- 
    phi_stmt_474_req_3518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_474_req_3518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(474), ack => phi_stmt_474_req_1); -- 
    convTranspose_cp_element_group_474: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_474"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(472) & convTranspose_CP_34_elements(473);
      gj_convTranspose_cp_element_group_474 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(474), clk => clk, reset => reset); --
    end block;
    -- CP-element group 475:  merge  transition  place  bypass 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	471 
    -- CP-element group 475: 	474 
    -- CP-element group 475: successors 
    -- CP-element group 475: 	476 
    -- CP-element group 475:  members (2) 
      -- CP-element group 475: 	 branch_block_stmt_38/merge_stmt_473_PhiReqMerge
      -- CP-element group 475: 	 branch_block_stmt_38/merge_stmt_473_PhiAck/$entry
      -- 
    convTranspose_CP_34_elements(475) <= OrReduce(convTranspose_CP_34_elements(471) & convTranspose_CP_34_elements(474));
    -- CP-element group 476:  fork  transition  place  input  output  bypass 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: 	475 
    -- CP-element group 476: successors 
    -- CP-element group 476: 	163 
    -- CP-element group 476: 	125 
    -- CP-element group 476: 	126 
    -- CP-element group 476: 	128 
    -- CP-element group 476: 	129 
    -- CP-element group 476: 	132 
    -- CP-element group 476: 	136 
    -- CP-element group 476: 	140 
    -- CP-element group 476: 	144 
    -- CP-element group 476: 	148 
    -- CP-element group 476: 	152 
    -- CP-element group 476: 	156 
    -- CP-element group 476: 	160 
    -- CP-element group 476:  members (56) 
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Update/cr
      -- CP-element group 476: 	 branch_block_stmt_38/merge_stmt_473__exit__
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636__entry__
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Update/cr
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_update_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_update_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/word_access_complete/word_0/cr
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/word_access_complete/word_0/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_update_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/word_access_complete/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Update/cr
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_update_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Update/cr
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_update_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_update_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Update/cr
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_update_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_resized_1
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_scaled_1
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_computed_1
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_resize_1/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_resize_1/$exit
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_resize_1/index_resize_req
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_resize_1/index_resize_ack
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_scale_1/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_scale_1/$exit
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_scale_1/scale_rename_req
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_scale_1/scale_rename_ack
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_update_start
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Sample/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Sample/req
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Update/req
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_complete/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_complete/req
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_sample_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Sample/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Sample/rr
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_update_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Update/cr
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_update_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Update/cr
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_update_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Update/cr
      -- CP-element group 476: 	 branch_block_stmt_38/merge_stmt_473_PhiAck/$exit
      -- CP-element group 476: 	 branch_block_stmt_38/merge_stmt_473_PhiAck/phi_stmt_474_ack
      -- 
    phi_stmt_474_ack_3523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 476_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_474_ack_0, ack => convTranspose_CP_34_elements(476)); -- 
    cr_1224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => type_cast_615_inst_req_1); -- 
    cr_1112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => type_cast_543_inst_req_1); -- 
    cr_1274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => ptr_deref_623_store_0_req_1); -- 
    cr_1168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => type_cast_579_inst_req_1); -- 
    cr_1140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => type_cast_561_inst_req_1); -- 
    cr_1196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => type_cast_597_inst_req_1); -- 
    req_980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => array_obj_ref_486_index_offset_req_0); -- 
    req_985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => array_obj_ref_486_index_offset_req_1); -- 
    req_1000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => addr_of_487_final_reg_req_1); -- 
    rr_1009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => RPIPE_ConvTranspose_input_pipe_490_inst_req_0); -- 
    cr_1028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => type_cast_494_inst_req_1); -- 
    cr_1056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => type_cast_507_inst_req_1); -- 
    cr_1084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => type_cast_525_inst_req_1); -- 
    -- CP-element group 477:  transition  output  delay-element  bypass 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	168 
    -- CP-element group 477: successors 
    -- CP-element group 477: 	481 
    -- CP-element group 477:  members (5) 
      -- CP-element group 477: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/$exit
      -- CP-element group 477: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_681/$exit
      -- CP-element group 477: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/$exit
      -- CP-element group 477: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_685_konst_delay_trans
      -- CP-element group 477: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_req
      -- 
    phi_stmt_681_req_3546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_681_req_3546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(477), ack => phi_stmt_681_req_0); -- 
    -- Element group convTranspose_CP_34_elements(477) is a control-delay.
    cp_element_477_delay: control_delay_element  generic map(name => " 477_delay", delay_value => 1)  port map(req => convTranspose_CP_34_elements(168), ack => convTranspose_CP_34_elements(477), clk => clk, reset =>reset);
    -- CP-element group 478:  transition  input  bypass 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: 	210 
    -- CP-element group 478: successors 
    -- CP-element group 478: 	480 
    -- CP-element group 478:  members (2) 
      -- CP-element group 478: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Sample/$exit
      -- CP-element group 478: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Sample/ra
      -- 
    ra_3566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 478_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_687_inst_ack_0, ack => convTranspose_CP_34_elements(478)); -- 
    -- CP-element group 479:  transition  input  bypass 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	210 
    -- CP-element group 479: successors 
    -- CP-element group 479: 	480 
    -- CP-element group 479:  members (2) 
      -- CP-element group 479: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Update/$exit
      -- CP-element group 479: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Update/ca
      -- 
    ca_3571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 479_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_687_inst_ack_1, ack => convTranspose_CP_34_elements(479)); -- 
    -- CP-element group 480:  join  transition  output  bypass 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: 	478 
    -- CP-element group 480: 	479 
    -- CP-element group 480: successors 
    -- CP-element group 480: 	481 
    -- CP-element group 480:  members (6) 
      -- CP-element group 480: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/$exit
      -- CP-element group 480: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/$exit
      -- CP-element group 480: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/$exit
      -- CP-element group 480: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/$exit
      -- CP-element group 480: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/$exit
      -- CP-element group 480: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_req
      -- 
    phi_stmt_681_req_3572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_681_req_3572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(480), ack => phi_stmt_681_req_1); -- 
    convTranspose_cp_element_group_480: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_480"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(478) & convTranspose_CP_34_elements(479);
      gj_convTranspose_cp_element_group_480 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(480), clk => clk, reset => reset); --
    end block;
    -- CP-element group 481:  merge  transition  place  bypass 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	477 
    -- CP-element group 481: 	480 
    -- CP-element group 481: successors 
    -- CP-element group 481: 	482 
    -- CP-element group 481:  members (2) 
      -- CP-element group 481: 	 branch_block_stmt_38/merge_stmt_680_PhiReqMerge
      -- CP-element group 481: 	 branch_block_stmt_38/merge_stmt_680_PhiAck/$entry
      -- 
    convTranspose_CP_34_elements(481) <= OrReduce(convTranspose_CP_34_elements(477) & convTranspose_CP_34_elements(480));
    -- CP-element group 482:  fork  transition  place  input  output  bypass 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	481 
    -- CP-element group 482: successors 
    -- CP-element group 482: 	196 
    -- CP-element group 482: 	200 
    -- CP-element group 482: 	204 
    -- CP-element group 482: 	207 
    -- CP-element group 482: 	188 
    -- CP-element group 482: 	192 
    -- CP-element group 482: 	169 
    -- CP-element group 482: 	170 
    -- CP-element group 482: 	172 
    -- CP-element group 482: 	173 
    -- CP-element group 482: 	176 
    -- CP-element group 482: 	180 
    -- CP-element group 482: 	184 
    -- CP-element group 482:  members (56) 
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/merge_stmt_680__exit__
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843__entry__
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Update/req
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Sample/req
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_update_start
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Sample/rr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_complete/req
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_scale_1/scale_rename_ack
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_complete/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_scale_1/scale_rename_req
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_sample_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_scale_1/$exit
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_scale_1/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_resize_1/index_resize_ack
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_resize_1/index_resize_req
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_resize_1/$exit
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_resize_1/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_computed_1
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_scaled_1
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_resized_1
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/word_access_complete/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/word_access_complete/word_0/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/word_access_complete/word_0/cr
      -- CP-element group 482: 	 branch_block_stmt_38/merge_stmt_680_PhiAck/$exit
      -- CP-element group 482: 	 branch_block_stmt_38/merge_stmt_680_PhiAck/phi_stmt_681_ack
      -- 
    phi_stmt_681_ack_3577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 482_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_681_ack_0, ack => convTranspose_CP_34_elements(482)); -- 
    req_1344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => array_obj_ref_693_index_offset_req_1); -- 
    req_1339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => array_obj_ref_693_index_offset_req_0); -- 
    cr_1415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_714_inst_req_1); -- 
    cr_1443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_732_inst_req_1); -- 
    rr_1368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => RPIPE_ConvTranspose_input_pipe_697_inst_req_0); -- 
    req_1359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => addr_of_694_final_reg_req_1); -- 
    cr_1387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_701_inst_req_1); -- 
    cr_1471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_750_inst_req_1); -- 
    cr_1499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_768_inst_req_1); -- 
    cr_1527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_786_inst_req_1); -- 
    cr_1555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_804_inst_req_1); -- 
    cr_1583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_822_inst_req_1); -- 
    cr_1633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => ptr_deref_830_store_0_req_1); -- 
    -- CP-element group 483:  merge  fork  transition  place  output  bypass 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: 	209 
    -- CP-element group 483: 	122 
    -- CP-element group 483: successors 
    -- CP-element group 483: 	211 
    -- CP-element group 483: 	212 
    -- CP-element group 483: 	213 
    -- CP-element group 483: 	214 
    -- CP-element group 483: 	215 
    -- CP-element group 483: 	216 
    -- CP-element group 483:  members (25) 
      -- CP-element group 483: 	 branch_block_stmt_38/merge_stmt_852__exit__
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880__entry__
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/$entry
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_sample_start_
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_update_start_
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Sample/$entry
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Sample/rr
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Update/$entry
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Update/cr
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_sample_start_
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_update_start_
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Sample/$entry
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Sample/rr
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Update/$entry
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Update/cr
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_sample_start_
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_update_start_
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Sample/$entry
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Sample/rr
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Update/$entry
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Update/cr
      -- CP-element group 483: 	 branch_block_stmt_38/merge_stmt_852_PhiReqMerge
      -- CP-element group 483: 	 branch_block_stmt_38/merge_stmt_852_PhiAck/$entry
      -- CP-element group 483: 	 branch_block_stmt_38/merge_stmt_852_PhiAck/$exit
      -- CP-element group 483: 	 branch_block_stmt_38/merge_stmt_852_PhiAck/dummy
      -- 
    rr_1664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(483), ack => type_cast_855_inst_req_0); -- 
    cr_1669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(483), ack => type_cast_855_inst_req_1); -- 
    rr_1678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(483), ack => type_cast_859_inst_req_0); -- 
    cr_1683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(483), ack => type_cast_859_inst_req_1); -- 
    rr_1692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(483), ack => type_cast_863_inst_req_0); -- 
    cr_1697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(483), ack => type_cast_863_inst_req_1); -- 
    convTranspose_CP_34_elements(483) <= OrReduce(convTranspose_CP_34_elements(209) & convTranspose_CP_34_elements(122));
    -- CP-element group 484:  transition  output  delay-element  bypass 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	221 
    -- CP-element group 484: successors 
    -- CP-element group 484: 	488 
    -- CP-element group 484:  members (5) 
      -- CP-element group 484: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/$exit
      -- CP-element group 484: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_925/$exit
      -- CP-element group 484: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/$exit
      -- CP-element group 484: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_931_konst_delay_trans
      -- CP-element group 484: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_req
      -- 
    phi_stmt_925_req_3623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_925_req_3623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(484), ack => phi_stmt_925_req_1); -- 
    -- Element group convTranspose_CP_34_elements(484) is a control-delay.
    cp_element_484_delay: control_delay_element  generic map(name => " 484_delay", delay_value => 1)  port map(req => convTranspose_CP_34_elements(221), ack => convTranspose_CP_34_elements(484), clk => clk, reset =>reset);
    -- CP-element group 485:  transition  input  bypass 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	230 
    -- CP-element group 485: successors 
    -- CP-element group 485: 	487 
    -- CP-element group 485:  members (2) 
      -- CP-element group 485: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Sample/$exit
      -- CP-element group 485: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Sample/ra
      -- 
    ra_3643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 485_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_928_inst_ack_0, ack => convTranspose_CP_34_elements(485)); -- 
    -- CP-element group 486:  transition  input  bypass 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: 	230 
    -- CP-element group 486: successors 
    -- CP-element group 486: 	487 
    -- CP-element group 486:  members (2) 
      -- CP-element group 486: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Update/$exit
      -- CP-element group 486: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Update/ca
      -- 
    ca_3648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 486_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_928_inst_ack_1, ack => convTranspose_CP_34_elements(486)); -- 
    -- CP-element group 487:  join  transition  output  bypass 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: 	485 
    -- CP-element group 487: 	486 
    -- CP-element group 487: successors 
    -- CP-element group 487: 	488 
    -- CP-element group 487:  members (6) 
      -- CP-element group 487: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/$exit
      -- CP-element group 487: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/$exit
      -- CP-element group 487: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/$exit
      -- CP-element group 487: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/$exit
      -- CP-element group 487: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/$exit
      -- CP-element group 487: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_req
      -- 
    phi_stmt_925_req_3649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_925_req_3649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(487), ack => phi_stmt_925_req_0); -- 
    convTranspose_cp_element_group_487: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_487"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(485) & convTranspose_CP_34_elements(486);
      gj_convTranspose_cp_element_group_487 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(487), clk => clk, reset => reset); --
    end block;
    -- CP-element group 488:  merge  transition  place  bypass 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: 	484 
    -- CP-element group 488: 	487 
    -- CP-element group 488: successors 
    -- CP-element group 488: 	489 
    -- CP-element group 488:  members (2) 
      -- CP-element group 488: 	 branch_block_stmt_38/merge_stmt_924_PhiReqMerge
      -- CP-element group 488: 	 branch_block_stmt_38/merge_stmt_924_PhiAck/$entry
      -- 
    convTranspose_CP_34_elements(488) <= OrReduce(convTranspose_CP_34_elements(484) & convTranspose_CP_34_elements(487));
    -- CP-element group 489:  fork  transition  place  input  output  bypass 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	488 
    -- CP-element group 489: successors 
    -- CP-element group 489: 	225 
    -- CP-element group 489: 	227 
    -- CP-element group 489: 	222 
    -- CP-element group 489: 	223 
    -- CP-element group 489:  members (29) 
      -- CP-element group 489: 	 branch_block_stmt_38/merge_stmt_924__exit__
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955__entry__
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_update_start_
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_resized_1
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_scaled_1
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_computed_1
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_resize_1/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_resize_1/$exit
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_resize_1/index_resize_req
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_resize_1/index_resize_ack
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_scale_1/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_scale_1/$exit
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_scale_1/scale_rename_req
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_scale_1/scale_rename_ack
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_update_start
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Sample/req
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Update/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Update/req
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_complete/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_complete/req
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_update_start_
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/word_access_complete/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/word_access_complete/word_0/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/word_access_complete/word_0/cr
      -- CP-element group 489: 	 branch_block_stmt_38/merge_stmt_924_PhiAck/$exit
      -- CP-element group 489: 	 branch_block_stmt_38/merge_stmt_924_PhiAck/phi_stmt_925_ack
      -- 
    phi_stmt_925_ack_3654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 489_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_925_ack_0, ack => convTranspose_CP_34_elements(489)); -- 
    req_1762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(489), ack => array_obj_ref_937_index_offset_req_0); -- 
    req_1767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(489), ack => array_obj_ref_937_index_offset_req_1); -- 
    req_1782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(489), ack => addr_of_938_final_reg_req_1); -- 
    cr_1832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(489), ack => ptr_deref_941_store_0_req_1); -- 
    -- CP-element group 490:  merge  fork  transition  place  output  bypass 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: 	229 
    -- CP-element group 490: 	219 
    -- CP-element group 490: successors 
    -- CP-element group 490: 	231 
    -- CP-element group 490: 	232 
    -- CP-element group 490: 	234 
    -- CP-element group 490:  members (16) 
      -- CP-element group 490: 	 branch_block_stmt_38/merge_stmt_964__exit__
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973__entry__
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/$entry
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_sample_start_
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_update_start_
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Sample/$entry
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Sample/crr
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Update/$entry
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Update/ccr
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_update_start_
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Update/$entry
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Update/cr
      -- CP-element group 490: 	 branch_block_stmt_38/merge_stmt_964_PhiReqMerge
      -- CP-element group 490: 	 branch_block_stmt_38/merge_stmt_964_PhiAck/$entry
      -- CP-element group 490: 	 branch_block_stmt_38/merge_stmt_964_PhiAck/$exit
      -- CP-element group 490: 	 branch_block_stmt_38/merge_stmt_964_PhiAck/dummy
      -- 
    crr_1863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(490), ack => call_stmt_967_call_req_0); -- 
    ccr_1868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(490), ack => call_stmt_967_call_req_1); -- 
    cr_1882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(490), ack => type_cast_972_inst_req_1); -- 
    convTranspose_CP_34_elements(490) <= OrReduce(convTranspose_CP_34_elements(229) & convTranspose_CP_34_elements(219));
    -- CP-element group 491:  transition  output  delay-element  bypass 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: 	421 
    -- CP-element group 491: successors 
    -- CP-element group 491: 	495 
    -- CP-element group 491:  members (5) 
      -- CP-element group 491: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/$exit
      -- CP-element group 491: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1356/$exit
      -- CP-element group 491: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/$exit
      -- CP-element group 491: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1360_konst_delay_trans
      -- CP-element group 491: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_req
      -- 
    phi_stmt_1356_req_3700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1356_req_3700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(491), ack => phi_stmt_1356_req_0); -- 
    -- Element group convTranspose_CP_34_elements(491) is a control-delay.
    cp_element_491_delay: control_delay_element  generic map(name => " 491_delay", delay_value => 1)  port map(req => convTranspose_CP_34_elements(421), ack => convTranspose_CP_34_elements(491), clk => clk, reset =>reset);
    -- CP-element group 492:  transition  input  bypass 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: 	469 
    -- CP-element group 492: successors 
    -- CP-element group 492: 	494 
    -- CP-element group 492:  members (2) 
      -- CP-element group 492: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/SplitProtocol/Sample/$exit
      -- CP-element group 492: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/SplitProtocol/Sample/ra
      -- 
    ra_3720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 492_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1362_inst_ack_0, ack => convTranspose_CP_34_elements(492)); -- 
    -- CP-element group 493:  transition  input  bypass 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	469 
    -- CP-element group 493: successors 
    -- CP-element group 493: 	494 
    -- CP-element group 493:  members (2) 
      -- CP-element group 493: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/SplitProtocol/Update/$exit
      -- CP-element group 493: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/SplitProtocol/Update/ca
      -- 
    ca_3725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 493_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1362_inst_ack_1, ack => convTranspose_CP_34_elements(493)); -- 
    -- CP-element group 494:  join  transition  output  bypass 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	492 
    -- CP-element group 494: 	493 
    -- CP-element group 494: successors 
    -- CP-element group 494: 	495 
    -- CP-element group 494:  members (6) 
      -- CP-element group 494: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/$exit
      -- CP-element group 494: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/$exit
      -- CP-element group 494: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/$exit
      -- CP-element group 494: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/$exit
      -- CP-element group 494: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/SplitProtocol/$exit
      -- CP-element group 494: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_req
      -- 
    phi_stmt_1356_req_3726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1356_req_3726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(494), ack => phi_stmt_1356_req_1); -- 
    convTranspose_cp_element_group_494: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_494"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(492) & convTranspose_CP_34_elements(493);
      gj_convTranspose_cp_element_group_494 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(494), clk => clk, reset => reset); --
    end block;
    -- CP-element group 495:  merge  transition  place  bypass 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	491 
    -- CP-element group 495: 	494 
    -- CP-element group 495: successors 
    -- CP-element group 495: 	496 
    -- CP-element group 495:  members (2) 
      -- CP-element group 495: 	 branch_block_stmt_38/merge_stmt_1355_PhiReqMerge
      -- CP-element group 495: 	 branch_block_stmt_38/merge_stmt_1355_PhiAck/$entry
      -- 
    convTranspose_CP_34_elements(495) <= OrReduce(convTranspose_CP_34_elements(491) & convTranspose_CP_34_elements(494));
    -- CP-element group 496:  fork  transition  place  input  output  bypass 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	495 
    -- CP-element group 496: successors 
    -- CP-element group 496: 	422 
    -- CP-element group 496: 	423 
    -- CP-element group 496: 	425 
    -- CP-element group 496: 	427 
    -- CP-element group 496: 	429 
    -- CP-element group 496: 	431 
    -- CP-element group 496: 	433 
    -- CP-element group 496: 	435 
    -- CP-element group 496: 	437 
    -- CP-element group 496: 	439 
    -- CP-element group 496: 	441 
    -- CP-element group 496: 	443 
    -- CP-element group 496:  members (53) 
      -- CP-element group 496: 	 branch_block_stmt_38/merge_stmt_1355__exit__
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483__entry__
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_update_start_
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/word_access_complete/word_0/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/word_access_complete/word_0/cr
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_Update/cr
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_scale_1/scale_rename_req
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_Update/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_update_start_
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_resize_1/index_resize_req
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_scale_1/$exit
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_Update/cr
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_resize_1/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/word_access_complete/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_update_start_
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_resized_1
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_Update/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_scaled_1
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_resize_1/$exit
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_resize_1/index_resize_ack
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_computed_1
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_update_start_
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_scale_1/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_scale_1/scale_rename_ack
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_Update/cr
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_update_start_
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_Update/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_Update/cr
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_Update/cr
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_Update/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_Update/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_update_start_
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_update_start_
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_update_start_
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_complete/req
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_complete/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_Update/cr
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_Update/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_Update/cr
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_update_start_
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_final_index_sum_regn_Update/req
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_update_start_
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_final_index_sum_regn_Update/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_Update/cr
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_Update/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_final_index_sum_regn_Sample/req
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_Update/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_final_index_sum_regn_Sample/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_final_index_sum_regn_update_start
      -- CP-element group 496: 	 branch_block_stmt_38/merge_stmt_1355_PhiAck/$exit
      -- CP-element group 496: 	 branch_block_stmt_38/merge_stmt_1355_PhiAck/phi_stmt_1356_ack
      -- 
    phi_stmt_1356_ack_3731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 496_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1356_ack_0, ack => convTranspose_CP_34_elements(496)); -- 
    cr_3197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => ptr_deref_1373_load_0_req_1); -- 
    cr_3272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => type_cast_1417_inst_req_1); -- 
    cr_3230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => type_cast_1387_inst_req_1); -- 
    cr_3286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => type_cast_1427_inst_req_1); -- 
    cr_3216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => type_cast_1377_inst_req_1); -- 
    cr_3258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => type_cast_1407_inst_req_1); -- 
    req_3152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => addr_of_1369_final_reg_req_1); -- 
    cr_3314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => type_cast_1447_inst_req_1); -- 
    cr_3244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => type_cast_1397_inst_req_1); -- 
    req_3137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => array_obj_ref_1368_index_offset_req_1); -- 
    cr_3300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => type_cast_1437_inst_req_1); -- 
    req_3132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => array_obj_ref_1368_index_offset_req_0); -- 
    -- CP-element group 497:  merge  transition  place  bypass 
    -- CP-element group 497: predecessors 
    -- CP-element group 497: 	419 
    -- CP-element group 497: 	468 
    -- CP-element group 497: successors 
    -- CP-element group 497:  members (16) 
      -- CP-element group 497: 	 $exit
      -- CP-element group 497: 	 branch_block_stmt_38/$exit
      -- CP-element group 497: 	 branch_block_stmt_38/branch_block_stmt_38__exit__
      -- CP-element group 497: 	 branch_block_stmt_38/merge_stmt_1492__exit__
      -- CP-element group 497: 	 branch_block_stmt_38/return__
      -- CP-element group 497: 	 branch_block_stmt_38/merge_stmt_1494__exit__
      -- CP-element group 497: 	 branch_block_stmt_38/merge_stmt_1492_PhiReqMerge
      -- CP-element group 497: 	 branch_block_stmt_38/merge_stmt_1492_PhiAck/$entry
      -- CP-element group 497: 	 branch_block_stmt_38/merge_stmt_1492_PhiAck/$exit
      -- CP-element group 497: 	 branch_block_stmt_38/merge_stmt_1492_PhiAck/dummy
      -- CP-element group 497: 	 branch_block_stmt_38/return___PhiReq/$entry
      -- CP-element group 497: 	 branch_block_stmt_38/return___PhiReq/$exit
      -- CP-element group 497: 	 branch_block_stmt_38/merge_stmt_1494_PhiReqMerge
      -- CP-element group 497: 	 branch_block_stmt_38/merge_stmt_1494_PhiAck/$entry
      -- CP-element group 497: 	 branch_block_stmt_38/merge_stmt_1494_PhiAck/$exit
      -- CP-element group 497: 	 branch_block_stmt_38/merge_stmt_1494_PhiAck/dummy
      -- 
    convTranspose_CP_34_elements(497) <= OrReduce(convTranspose_CP_34_elements(419) & convTranspose_CP_34_elements(468));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar525_936_resized : std_logic_vector(13 downto 0);
    signal R_indvar525_936_scaled : std_logic_vector(13 downto 0);
    signal R_indvar539_692_resized : std_logic_vector(10 downto 0);
    signal R_indvar539_692_scaled : std_logic_vector(10 downto 0);
    signal R_indvar555_485_resized : std_logic_vector(13 downto 0);
    signal R_indvar555_485_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1367_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1367_scaled : std_logic_vector(13 downto 0);
    signal add108_339 : std_logic_vector(15 downto 0);
    signal add117_364 : std_logic_vector(15 downto 0);
    signal add126_389 : std_logic_vector(15 downto 0);
    signal add12_88 : std_logic_vector(15 downto 0);
    signal add135_414 : std_logic_vector(15 downto 0);
    signal add150_513 : std_logic_vector(63 downto 0);
    signal add156_531 : std_logic_vector(63 downto 0);
    signal add162_549 : std_logic_vector(63 downto 0);
    signal add168_567 : std_logic_vector(63 downto 0);
    signal add174_585 : std_logic_vector(63 downto 0);
    signal add180_603 : std_logic_vector(63 downto 0);
    signal add186_621 : std_logic_vector(63 downto 0);
    signal add206_720 : std_logic_vector(63 downto 0);
    signal add212_738 : std_logic_vector(63 downto 0);
    signal add218_756 : std_logic_vector(63 downto 0);
    signal add21_113 : std_logic_vector(15 downto 0);
    signal add224_774 : std_logic_vector(63 downto 0);
    signal add230_792 : std_logic_vector(63 downto 0);
    signal add236_810 : std_logic_vector(63 downto 0);
    signal add242_828 : std_logic_vector(63 downto 0);
    signal add30_138 : std_logic_vector(15 downto 0);
    signal add39_163 : std_logic_vector(15 downto 0);
    signal add48_188 : std_logic_vector(15 downto 0);
    signal add57_213 : std_logic_vector(15 downto 0);
    signal add74_253 : std_logic_vector(31 downto 0);
    signal add79_258 : std_logic_vector(31 downto 0);
    signal add99_314 : std_logic_vector(15 downto 0);
    signal add_63 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1368_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1368_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1368_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1368_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1368_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1368_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_486_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_486_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_486_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_486_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_486_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_486_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_693_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_693_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_693_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_693_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_693_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_693_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_937_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_937_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_937_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_937_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_937_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_937_root_address : std_logic_vector(13 downto 0);
    signal arrayidx246_695 : std_logic_vector(31 downto 0);
    signal arrayidx269_939 : std_logic_vector(31 downto 0);
    signal arrayidx432_1370 : std_logic_vector(31 downto 0);
    signal arrayidx_488 : std_logic_vector(31 downto 0);
    signal call101_317 : std_logic_vector(7 downto 0);
    signal call106_330 : std_logic_vector(7 downto 0);
    signal call10_79 : std_logic_vector(7 downto 0);
    signal call110_342 : std_logic_vector(7 downto 0);
    signal call115_355 : std_logic_vector(7 downto 0);
    signal call119_367 : std_logic_vector(7 downto 0);
    signal call124_380 : std_logic_vector(7 downto 0);
    signal call128_392 : std_logic_vector(7 downto 0);
    signal call133_405 : std_logic_vector(7 downto 0);
    signal call143_491 : std_logic_vector(7 downto 0);
    signal call147_504 : std_logic_vector(7 downto 0);
    signal call14_91 : std_logic_vector(7 downto 0);
    signal call153_522 : std_logic_vector(7 downto 0);
    signal call159_540 : std_logic_vector(7 downto 0);
    signal call165_558 : std_logic_vector(7 downto 0);
    signal call171_576 : std_logic_vector(7 downto 0);
    signal call177_594 : std_logic_vector(7 downto 0);
    signal call183_612 : std_logic_vector(7 downto 0);
    signal call199_698 : std_logic_vector(7 downto 0);
    signal call19_104 : std_logic_vector(7 downto 0);
    signal call203_711 : std_logic_vector(7 downto 0);
    signal call209_729 : std_logic_vector(7 downto 0);
    signal call215_747 : std_logic_vector(7 downto 0);
    signal call221_765 : std_logic_vector(7 downto 0);
    signal call227_783 : std_logic_vector(7 downto 0);
    signal call233_801 : std_logic_vector(7 downto 0);
    signal call239_819 : std_logic_vector(7 downto 0);
    signal call23_116 : std_logic_vector(7 downto 0);
    signal call275_967 : std_logic_vector(63 downto 0);
    signal call28_129 : std_logic_vector(7 downto 0);
    signal call2_54 : std_logic_vector(7 downto 0);
    signal call32_141 : std_logic_vector(7 downto 0);
    signal call346_1190 : std_logic_vector(15 downto 0);
    signal call348_1193 : std_logic_vector(15 downto 0);
    signal call350_1196 : std_logic_vector(15 downto 0);
    signal call352_1199 : std_logic_vector(15 downto 0);
    signal call354_1202 : std_logic_vector(63 downto 0);
    signal call37_154 : std_logic_vector(7 downto 0);
    signal call41_166 : std_logic_vector(7 downto 0);
    signal call46_179 : std_logic_vector(7 downto 0);
    signal call50_191 : std_logic_vector(7 downto 0);
    signal call55_204 : std_logic_vector(7 downto 0);
    signal call5_66 : std_logic_vector(7 downto 0);
    signal call92_292 : std_logic_vector(7 downto 0);
    signal call97_305 : std_logic_vector(7 downto 0);
    signal call_41 : std_logic_vector(7 downto 0);
    signal cmp194509_435 : std_logic_vector(0 downto 0);
    signal cmp264505_880 : std_logic_vector(0 downto 0);
    signal cmp513_420 : std_logic_vector(0 downto 0);
    signal conv104_321 : std_logic_vector(15 downto 0);
    signal conv107_334 : std_logic_vector(15 downto 0);
    signal conv113_346 : std_logic_vector(15 downto 0);
    signal conv116_359 : std_logic_vector(15 downto 0);
    signal conv11_83 : std_logic_vector(15 downto 0);
    signal conv122_371 : std_logic_vector(15 downto 0);
    signal conv125_384 : std_logic_vector(15 downto 0);
    signal conv131_396 : std_logic_vector(15 downto 0);
    signal conv134_409 : std_logic_vector(15 downto 0);
    signal conv144_495 : std_logic_vector(63 downto 0);
    signal conv149_508 : std_logic_vector(63 downto 0);
    signal conv155_526 : std_logic_vector(63 downto 0);
    signal conv161_544 : std_logic_vector(63 downto 0);
    signal conv167_562 : std_logic_vector(63 downto 0);
    signal conv173_580 : std_logic_vector(63 downto 0);
    signal conv179_598 : std_logic_vector(63 downto 0);
    signal conv17_95 : std_logic_vector(15 downto 0);
    signal conv185_616 : std_logic_vector(63 downto 0);
    signal conv1_45 : std_logic_vector(15 downto 0);
    signal conv200_702 : std_logic_vector(63 downto 0);
    signal conv205_715 : std_logic_vector(63 downto 0);
    signal conv20_108 : std_logic_vector(15 downto 0);
    signal conv211_733 : std_logic_vector(63 downto 0);
    signal conv217_751 : std_logic_vector(63 downto 0);
    signal conv223_769 : std_logic_vector(63 downto 0);
    signal conv229_787 : std_logic_vector(63 downto 0);
    signal conv235_805 : std_logic_vector(63 downto 0);
    signal conv241_823 : std_logic_vector(63 downto 0);
    signal conv253_856 : std_logic_vector(31 downto 0);
    signal conv255_860 : std_logic_vector(31 downto 0);
    signal conv258_864 : std_logic_vector(31 downto 0);
    signal conv26_120 : std_logic_vector(15 downto 0);
    signal conv276_973 : std_logic_vector(63 downto 0);
    signal conv29_133 : std_logic_vector(15 downto 0);
    signal conv305_1055 : std_logic_vector(15 downto 0);
    signal conv307_1062 : std_logic_vector(15 downto 0);
    signal conv322_1111 : std_logic_vector(15 downto 0);
    signal conv324_1118 : std_logic_vector(15 downto 0);
    signal conv339_1167 : std_logic_vector(15 downto 0);
    signal conv341_1174 : std_logic_vector(15 downto 0);
    signal conv355_1207 : std_logic_vector(63 downto 0);
    signal conv35_145 : std_logic_vector(15 downto 0);
    signal conv361_1216 : std_logic_vector(7 downto 0);
    signal conv367_1226 : std_logic_vector(7 downto 0);
    signal conv373_1236 : std_logic_vector(7 downto 0);
    signal conv379_1246 : std_logic_vector(7 downto 0);
    signal conv385_1256 : std_logic_vector(7 downto 0);
    signal conv38_158 : std_logic_vector(15 downto 0);
    signal conv391_1266 : std_logic_vector(7 downto 0);
    signal conv397_1276 : std_logic_vector(7 downto 0);
    signal conv3_58 : std_logic_vector(15 downto 0);
    signal conv403_1286 : std_logic_vector(7 downto 0);
    signal conv437_1378 : std_logic_vector(7 downto 0);
    signal conv443_1388 : std_logic_vector(7 downto 0);
    signal conv449_1398 : std_logic_vector(7 downto 0);
    signal conv44_170 : std_logic_vector(15 downto 0);
    signal conv455_1408 : std_logic_vector(7 downto 0);
    signal conv461_1418 : std_logic_vector(7 downto 0);
    signal conv467_1428 : std_logic_vector(7 downto 0);
    signal conv473_1438 : std_logic_vector(7 downto 0);
    signal conv479_1448 : std_logic_vector(7 downto 0);
    signal conv47_183 : std_logic_vector(15 downto 0);
    signal conv53_195 : std_logic_vector(15 downto 0);
    signal conv56_208 : std_logic_vector(15 downto 0);
    signal conv61_217 : std_logic_vector(31 downto 0);
    signal conv63_221 : std_logic_vector(31 downto 0);
    signal conv65_225 : std_logic_vector(31 downto 0);
    signal conv82_262 : std_logic_vector(31 downto 0);
    signal conv84_266 : std_logic_vector(31 downto 0);
    signal conv87_270 : std_logic_vector(31 downto 0);
    signal conv8_70 : std_logic_vector(15 downto 0);
    signal conv90_274 : std_logic_vector(31 downto 0);
    signal conv95_296 : std_logic_vector(15 downto 0);
    signal conv98_309 : std_logic_vector(15 downto 0);
    signal exitcond1_1483 : std_logic_vector(0 downto 0);
    signal exitcond2_843 : std_logic_vector(0 downto 0);
    signal exitcond3_636 : std_logic_vector(0 downto 0);
    signal exitcond_955 : std_logic_vector(0 downto 0);
    signal iNsTr_14_247 : std_logic_vector(31 downto 0);
    signal iNsTr_196_1340 : std_logic_vector(63 downto 0);
    signal iNsTr_26_458 : std_logic_vector(63 downto 0);
    signal iNsTr_39_665 : std_logic_vector(63 downto 0);
    signal iNsTr_53_909 : std_logic_vector(63 downto 0);
    signal indvar525_925 : std_logic_vector(63 downto 0);
    signal indvar539_681 : std_logic_vector(63 downto 0);
    signal indvar555_474 : std_logic_vector(63 downto 0);
    signal indvar_1356 : std_logic_vector(63 downto 0);
    signal indvarx_xnext526_950 : std_logic_vector(63 downto 0);
    signal indvarx_xnext540_838 : std_logic_vector(63 downto 0);
    signal indvarx_xnext556_631 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1478 : std_logic_vector(63 downto 0);
    signal mul256_869 : std_logic_vector(31 downto 0);
    signal mul259_874 : std_logic_vector(31 downto 0);
    signal mul66_235 : std_logic_vector(31 downto 0);
    signal mul85_279 : std_logic_vector(31 downto 0);
    signal mul88_284 : std_logic_vector(31 downto 0);
    signal mul91_289 : std_logic_vector(31 downto 0);
    signal mul_230 : std_logic_vector(31 downto 0);
    signal ptr_deref_1373_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1373_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1373_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1373_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1373_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_623_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_623_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_623_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_623_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_623_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_623_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_830_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_830_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_830_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_830_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_830_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_830_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_941_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_941_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_941_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_941_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_941_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_941_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl105_327 : std_logic_vector(15 downto 0);
    signal shl114_352 : std_logic_vector(15 downto 0);
    signal shl123_377 : std_logic_vector(15 downto 0);
    signal shl132_402 : std_logic_vector(15 downto 0);
    signal shl146_501 : std_logic_vector(63 downto 0);
    signal shl152_519 : std_logic_vector(63 downto 0);
    signal shl158_537 : std_logic_vector(63 downto 0);
    signal shl164_555 : std_logic_vector(63 downto 0);
    signal shl170_573 : std_logic_vector(63 downto 0);
    signal shl176_591 : std_logic_vector(63 downto 0);
    signal shl182_609 : std_logic_vector(63 downto 0);
    signal shl18_101 : std_logic_vector(15 downto 0);
    signal shl202_708 : std_logic_vector(63 downto 0);
    signal shl208_726 : std_logic_vector(63 downto 0);
    signal shl214_744 : std_logic_vector(63 downto 0);
    signal shl220_762 : std_logic_vector(63 downto 0);
    signal shl226_780 : std_logic_vector(63 downto 0);
    signal shl232_798 : std_logic_vector(63 downto 0);
    signal shl238_816 : std_logic_vector(63 downto 0);
    signal shl27_126 : std_logic_vector(15 downto 0);
    signal shl36_151 : std_logic_vector(15 downto 0);
    signal shl45_176 : std_logic_vector(15 downto 0);
    signal shl54_201 : std_logic_vector(15 downto 0);
    signal shl96_302 : std_logic_vector(15 downto 0);
    signal shl9_76 : std_logic_vector(15 downto 0);
    signal shl_51 : std_logic_vector(15 downto 0);
    signal shr304_1051 : std_logic_vector(31 downto 0);
    signal shr321_1107 : std_logic_vector(31 downto 0);
    signal shr338_1163 : std_logic_vector(31 downto 0);
    signal shr364_1222 : std_logic_vector(63 downto 0);
    signal shr370_1232 : std_logic_vector(63 downto 0);
    signal shr376_1242 : std_logic_vector(63 downto 0);
    signal shr382_1252 : std_logic_vector(63 downto 0);
    signal shr388_1262 : std_logic_vector(63 downto 0);
    signal shr394_1272 : std_logic_vector(63 downto 0);
    signal shr400_1282 : std_logic_vector(63 downto 0);
    signal shr440_1384 : std_logic_vector(63 downto 0);
    signal shr446_1394 : std_logic_vector(63 downto 0);
    signal shr452_1404 : std_logic_vector(63 downto 0);
    signal shr458_1414 : std_logic_vector(63 downto 0);
    signal shr464_1424 : std_logic_vector(63 downto 0);
    signal shr470_1434 : std_logic_vector(63 downto 0);
    signal shr476_1444 : std_logic_vector(63 downto 0);
    signal shr_241 : std_logic_vector(31 downto 0);
    signal sub_1212 : std_logic_vector(63 downto 0);
    signal tmp433_1374 : std_logic_vector(63 downto 0);
    signal tmp520_1324 : std_logic_vector(31 downto 0);
    signal tmp520x_xop_1336 : std_logic_vector(31 downto 0);
    signal tmp521_1330 : std_logic_vector(0 downto 0);
    signal tmp524_1353 : std_logic_vector(63 downto 0);
    signal tmp532_893 : std_logic_vector(31 downto 0);
    signal tmp532x_xop_905 : std_logic_vector(31 downto 0);
    signal tmp533_899 : std_logic_vector(0 downto 0);
    signal tmp537_922 : std_logic_vector(63 downto 0);
    signal tmp548_649 : std_logic_vector(31 downto 0);
    signal tmp548x_xop_661 : std_logic_vector(31 downto 0);
    signal tmp549_655 : std_logic_vector(0 downto 0);
    signal tmp553_678 : std_logic_vector(63 downto 0);
    signal tmp562x_xop_454 : std_logic_vector(31 downto 0);
    signal tmp563_448 : std_logic_vector(0 downto 0);
    signal tmp567_471 : std_logic_vector(63 downto 0);
    signal type_cast_1004_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1008_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1049_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1105_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1161_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1205_wire : std_logic_vector(63 downto 0);
    signal type_cast_1220_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1230_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1240_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_124_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1250_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1260_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1270_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1280_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1322_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1328_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1334_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1344_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1351_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1360_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1362_wire : std_logic_vector(63 downto 0);
    signal type_cast_1382_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1392_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1402_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1412_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1422_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1432_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1442_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1476_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_149_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_174_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_199_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_239_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_245_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_251_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_300_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_325_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_350_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_375_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_400_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_418_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_433_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_446_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_452_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_462_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_469_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_478_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_480_wire : std_logic_vector(63 downto 0);
    signal type_cast_499_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_49_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_517_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_535_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_553_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_571_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_589_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_607_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_629_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_647_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_653_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_659_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_669_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_676_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_685_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_687_wire : std_logic_vector(63 downto 0);
    signal type_cast_706_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_724_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_742_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_74_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_760_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_778_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_796_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_814_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_836_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_878_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_891_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_897_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_903_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_913_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_920_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_928_wire : std_logic_vector(63 downto 0);
    signal type_cast_931_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_943_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_948_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_971_wire : std_logic_vector(63 downto 0);
    signal type_cast_99_wire_constant : std_logic_vector(15 downto 0);
    signal xx_xop569_915 : std_logic_vector(63 downto 0);
    signal xx_xop570_671 : std_logic_vector(63 downto 0);
    signal xx_xop571_464 : std_logic_vector(63 downto 0);
    signal xx_xop_1346 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1368_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1368_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1368_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1368_resized_base_address <= "00000000000000";
    array_obj_ref_486_constant_part_of_offset <= "00000000000000";
    array_obj_ref_486_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_486_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_486_resized_base_address <= "00000000000000";
    array_obj_ref_693_constant_part_of_offset <= "00000100010";
    array_obj_ref_693_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_693_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_693_resized_base_address <= "00000000000";
    array_obj_ref_937_constant_part_of_offset <= "00000000000000";
    array_obj_ref_937_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_937_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_937_resized_base_address <= "00000000000000";
    ptr_deref_1373_word_offset_0 <= "00000000000000";
    ptr_deref_623_word_offset_0 <= "00000000000000";
    ptr_deref_830_word_offset_0 <= "00000000000";
    ptr_deref_941_word_offset_0 <= "00000000000000";
    type_cast_1004_wire_constant <= "0000000000000000";
    type_cast_1008_wire_constant <= "0000000000000000";
    type_cast_1049_wire_constant <= "00000000000000000000000000010010";
    type_cast_1105_wire_constant <= "00000000000000000000000000010001";
    type_cast_1161_wire_constant <= "00000000000000000000000000010000";
    type_cast_1220_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1230_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1240_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_124_wire_constant <= "0000000000001000";
    type_cast_1250_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1260_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1270_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1280_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1322_wire_constant <= "00000000000000000000000000000010";
    type_cast_1328_wire_constant <= "00000000000000000000000000000001";
    type_cast_1334_wire_constant <= "11111111111111111111111111111111";
    type_cast_1344_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1351_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1360_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1382_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1392_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1402_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1412_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1422_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1432_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1442_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1476_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_149_wire_constant <= "0000000000001000";
    type_cast_174_wire_constant <= "0000000000001000";
    type_cast_199_wire_constant <= "0000000000001000";
    type_cast_239_wire_constant <= "00000000000000000000000000000010";
    type_cast_245_wire_constant <= "00000000000000000000000000000001";
    type_cast_251_wire_constant <= "01111111111111111111111111111110";
    type_cast_300_wire_constant <= "0000000000001000";
    type_cast_325_wire_constant <= "0000000000001000";
    type_cast_350_wire_constant <= "0000000000001000";
    type_cast_375_wire_constant <= "0000000000001000";
    type_cast_400_wire_constant <= "0000000000001000";
    type_cast_418_wire_constant <= "00000000000000000000000000000011";
    type_cast_433_wire_constant <= "00000000000000000000000000000011";
    type_cast_446_wire_constant <= "00000000000000000000000000000001";
    type_cast_452_wire_constant <= "11111111111111111111111111111111";
    type_cast_462_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_469_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_478_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_499_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_49_wire_constant <= "0000000000001000";
    type_cast_517_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_535_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_553_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_571_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_589_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_607_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_629_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_647_wire_constant <= "00000000000000000000000000000010";
    type_cast_653_wire_constant <= "00000000000000000000000000000001";
    type_cast_659_wire_constant <= "11111111111111111111111111111111";
    type_cast_669_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_676_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_685_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_706_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_724_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_742_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_74_wire_constant <= "0000000000001000";
    type_cast_760_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_778_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_796_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_814_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_836_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_878_wire_constant <= "00000000000000000000000000000011";
    type_cast_891_wire_constant <= "00000000000000000000000000000010";
    type_cast_897_wire_constant <= "00000000000000000000000000000001";
    type_cast_903_wire_constant <= "11111111111111111111111111111111";
    type_cast_913_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_920_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_931_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_943_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_948_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_99_wire_constant <= "0000000000001000";
    phi_stmt_1356: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1360_wire_constant & type_cast_1362_wire;
      req <= phi_stmt_1356_req_0 & phi_stmt_1356_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1356",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1356_ack_0,
          idata => idata,
          odata => indvar_1356,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1356
    phi_stmt_474: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_478_wire_constant & type_cast_480_wire;
      req <= phi_stmt_474_req_0 & phi_stmt_474_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_474",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_474_ack_0,
          idata => idata,
          odata => indvar555_474,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_474
    phi_stmt_681: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_685_wire_constant & type_cast_687_wire;
      req <= phi_stmt_681_req_0 & phi_stmt_681_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_681",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_681_ack_0,
          idata => idata,
          odata => indvar539_681,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_681
    phi_stmt_925: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_928_wire & type_cast_931_wire_constant;
      req <= phi_stmt_925_req_0 & phi_stmt_925_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_925",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_925_ack_0,
          idata => idata,
          odata => indvar525_925,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_925
    -- flow-through select operator MUX_1352_inst
    tmp524_1353 <= xx_xop_1346 when (tmp521_1330(0) /=  '0') else type_cast_1351_wire_constant;
    -- flow-through select operator MUX_470_inst
    tmp567_471 <= xx_xop571_464 when (tmp563_448(0) /=  '0') else type_cast_469_wire_constant;
    -- flow-through select operator MUX_677_inst
    tmp553_678 <= xx_xop570_671 when (tmp549_655(0) /=  '0') else type_cast_676_wire_constant;
    -- flow-through select operator MUX_921_inst
    tmp537_922 <= xx_xop569_915 when (tmp533_899(0) /=  '0') else type_cast_920_wire_constant;
    addr_of_1369_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1369_final_reg_req_0;
      addr_of_1369_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1369_final_reg_req_1;
      addr_of_1369_final_reg_ack_1<= rack(0);
      addr_of_1369_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1369_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1368_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx432_1370,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_487_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_487_final_reg_req_0;
      addr_of_487_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_487_final_reg_req_1;
      addr_of_487_final_reg_ack_1<= rack(0);
      addr_of_487_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_487_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_486_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_488,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_694_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_694_final_reg_req_0;
      addr_of_694_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_694_final_reg_req_1;
      addr_of_694_final_reg_ack_1<= rack(0);
      addr_of_694_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_694_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_693_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx246_695,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_938_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_938_final_reg_req_0;
      addr_of_938_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_938_final_reg_req_1;
      addr_of_938_final_reg_ack_1<= rack(0);
      addr_of_938_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_938_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_937_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx269_939,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1054_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1054_inst_req_0;
      type_cast_1054_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1054_inst_req_1;
      type_cast_1054_inst_ack_1<= rack(0);
      type_cast_1054_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1054_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr304_1051,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv305_1055,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1061_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1061_inst_req_0;
      type_cast_1061_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1061_inst_req_1;
      type_cast_1061_inst_ack_1<= rack(0);
      type_cast_1061_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1061_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_241,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv307_1062,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_107_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_107_inst_req_0;
      type_cast_107_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_107_inst_req_1;
      type_cast_107_inst_ack_1<= rack(0);
      type_cast_107_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_107_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_104,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_108,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1110_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1110_inst_req_0;
      type_cast_1110_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1110_inst_req_1;
      type_cast_1110_inst_ack_1<= rack(0);
      type_cast_1110_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1110_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr321_1107,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv322_1111,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1117_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1117_inst_req_0;
      type_cast_1117_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1117_inst_req_1;
      type_cast_1117_inst_ack_1<= rack(0);
      type_cast_1117_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1117_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add74_253,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv324_1118,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1166_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1166_inst_req_0;
      type_cast_1166_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1166_inst_req_1;
      type_cast_1166_inst_ack_1<= rack(0);
      type_cast_1166_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1166_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr338_1163,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv339_1167,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1173_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1173_inst_req_0;
      type_cast_1173_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1173_inst_req_1;
      type_cast_1173_inst_ack_1<= rack(0);
      type_cast_1173_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1173_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add79_258,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv341_1174,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_119_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_119_inst_req_0;
      type_cast_119_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_119_inst_req_1;
      type_cast_119_inst_ack_1<= rack(0);
      type_cast_119_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_119_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_116,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_120,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1206_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1206_inst_req_0;
      type_cast_1206_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1206_inst_req_1;
      type_cast_1206_inst_ack_1<= rack(0);
      type_cast_1206_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1206_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1205_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv355_1207,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1215_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1215_inst_req_0;
      type_cast_1215_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1215_inst_req_1;
      type_cast_1215_inst_ack_1<= rack(0);
      type_cast_1215_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1215_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_1212,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv361_1216,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1225_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1225_inst_req_0;
      type_cast_1225_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1225_inst_req_1;
      type_cast_1225_inst_ack_1<= rack(0);
      type_cast_1225_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1225_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr364_1222,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv367_1226,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1235_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1235_inst_req_0;
      type_cast_1235_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1235_inst_req_1;
      type_cast_1235_inst_ack_1<= rack(0);
      type_cast_1235_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1235_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr370_1232,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv373_1236,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1245_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1245_inst_req_0;
      type_cast_1245_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1245_inst_req_1;
      type_cast_1245_inst_ack_1<= rack(0);
      type_cast_1245_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1245_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr376_1242,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv379_1246,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1255_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1255_inst_req_0;
      type_cast_1255_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1255_inst_req_1;
      type_cast_1255_inst_ack_1<= rack(0);
      type_cast_1255_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1255_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr382_1252,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv385_1256,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1265_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1265_inst_req_0;
      type_cast_1265_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1265_inst_req_1;
      type_cast_1265_inst_ack_1<= rack(0);
      type_cast_1265_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1265_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr388_1262,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv391_1266,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1275_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1275_inst_req_0;
      type_cast_1275_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1275_inst_req_1;
      type_cast_1275_inst_ack_1<= rack(0);
      type_cast_1275_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1275_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr394_1272,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv397_1276,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1285_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1285_inst_req_0;
      type_cast_1285_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1285_inst_req_1;
      type_cast_1285_inst_ack_1<= rack(0);
      type_cast_1285_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1285_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr400_1282,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv403_1286,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_132_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_132_inst_req_0;
      type_cast_132_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_132_inst_req_1;
      type_cast_132_inst_ack_1<= rack(0);
      type_cast_132_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_132_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_129,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_133,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1339_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1339_inst_req_0;
      type_cast_1339_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1339_inst_req_1;
      type_cast_1339_inst_ack_1<= rack(0);
      type_cast_1339_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1339_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp520x_xop_1336,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_196_1340,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1362_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1362_inst_req_0;
      type_cast_1362_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1362_inst_req_1;
      type_cast_1362_inst_ack_1<= rack(0);
      type_cast_1362_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1362_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1478,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1362_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1377_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1377_inst_req_0;
      type_cast_1377_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1377_inst_req_1;
      type_cast_1377_inst_ack_1<= rack(0);
      type_cast_1377_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1377_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp433_1374,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv437_1378,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1387_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1387_inst_req_0;
      type_cast_1387_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1387_inst_req_1;
      type_cast_1387_inst_ack_1<= rack(0);
      type_cast_1387_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1387_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr440_1384,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv443_1388,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1397_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1397_inst_req_0;
      type_cast_1397_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1397_inst_req_1;
      type_cast_1397_inst_ack_1<= rack(0);
      type_cast_1397_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1397_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr446_1394,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv449_1398,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1407_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1407_inst_req_0;
      type_cast_1407_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1407_inst_req_1;
      type_cast_1407_inst_ack_1<= rack(0);
      type_cast_1407_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1407_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr452_1404,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv455_1408,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1417_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1417_inst_req_0;
      type_cast_1417_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1417_inst_req_1;
      type_cast_1417_inst_ack_1<= rack(0);
      type_cast_1417_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1417_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr458_1414,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv461_1418,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1427_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1427_inst_req_0;
      type_cast_1427_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1427_inst_req_1;
      type_cast_1427_inst_ack_1<= rack(0);
      type_cast_1427_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1427_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr464_1424,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv467_1428,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1437_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1437_inst_req_0;
      type_cast_1437_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1437_inst_req_1;
      type_cast_1437_inst_ack_1<= rack(0);
      type_cast_1437_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1437_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr470_1434,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv473_1438,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1447_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1447_inst_req_0;
      type_cast_1447_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1447_inst_req_1;
      type_cast_1447_inst_ack_1<= rack(0);
      type_cast_1447_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1447_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr476_1444,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv479_1448,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_144_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_144_inst_req_0;
      type_cast_144_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_144_inst_req_1;
      type_cast_144_inst_ack_1<= rack(0);
      type_cast_144_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_144_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_141,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_145,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_157_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_157_inst_req_0;
      type_cast_157_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_157_inst_req_1;
      type_cast_157_inst_ack_1<= rack(0);
      type_cast_157_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_157_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_154,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_158,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_169_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_169_inst_req_0;
      type_cast_169_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_169_inst_req_1;
      type_cast_169_inst_ack_1<= rack(0);
      type_cast_169_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_169_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_166,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_170,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_182_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_182_inst_req_0;
      type_cast_182_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_182_inst_req_1;
      type_cast_182_inst_ack_1<= rack(0);
      type_cast_182_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_182_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_179,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_183,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_194_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_194_inst_req_0;
      type_cast_194_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_194_inst_req_1;
      type_cast_194_inst_ack_1<= rack(0);
      type_cast_194_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_194_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_191,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_195,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_207_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_207_inst_req_0;
      type_cast_207_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_207_inst_req_1;
      type_cast_207_inst_ack_1<= rack(0);
      type_cast_207_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_207_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_204,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_208,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_216_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_216_inst_req_0;
      type_cast_216_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_216_inst_req_1;
      type_cast_216_inst_ack_1<= rack(0);
      type_cast_216_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_216_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_63,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_217,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_220_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_220_inst_req_0;
      type_cast_220_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_220_inst_req_1;
      type_cast_220_inst_ack_1<= rack(0);
      type_cast_220_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_220_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add12_88,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_221,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_224_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_224_inst_req_0;
      type_cast_224_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_224_inst_req_1;
      type_cast_224_inst_ack_1<= rack(0);
      type_cast_224_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_224_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_113,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_225,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_261_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_261_inst_req_0;
      type_cast_261_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_261_inst_req_1;
      type_cast_261_inst_ack_1<= rack(0);
      type_cast_261_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_261_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add30_138,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_262,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_265_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_265_inst_req_0;
      type_cast_265_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_265_inst_req_1;
      type_cast_265_inst_ack_1<= rack(0);
      type_cast_265_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_265_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add39_163,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_266,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_269_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_269_inst_req_0;
      type_cast_269_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_269_inst_req_1;
      type_cast_269_inst_ack_1<= rack(0);
      type_cast_269_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_269_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add48_188,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv87_270,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_273_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_273_inst_req_0;
      type_cast_273_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_273_inst_req_1;
      type_cast_273_inst_ack_1<= rack(0);
      type_cast_273_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_273_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add57_213,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_274,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_295_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_295_inst_req_0;
      type_cast_295_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_295_inst_req_1;
      type_cast_295_inst_ack_1<= rack(0);
      type_cast_295_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_295_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call92_292,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_296,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_308_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_308_inst_req_0;
      type_cast_308_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_308_inst_req_1;
      type_cast_308_inst_ack_1<= rack(0);
      type_cast_308_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_308_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_305,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_309,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_320_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_320_inst_req_0;
      type_cast_320_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_320_inst_req_1;
      type_cast_320_inst_ack_1<= rack(0);
      type_cast_320_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_320_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_317,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_321,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_333_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_333_inst_req_0;
      type_cast_333_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_333_inst_req_1;
      type_cast_333_inst_ack_1<= rack(0);
      type_cast_333_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_333_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_330,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_334,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_345_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_345_inst_req_0;
      type_cast_345_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_345_inst_req_1;
      type_cast_345_inst_ack_1<= rack(0);
      type_cast_345_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_345_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call110_342,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_346,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_358_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_358_inst_req_0;
      type_cast_358_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_358_inst_req_1;
      type_cast_358_inst_ack_1<= rack(0);
      type_cast_358_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_358_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_355,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_359,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_370_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_370_inst_req_0;
      type_cast_370_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_370_inst_req_1;
      type_cast_370_inst_ack_1<= rack(0);
      type_cast_370_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_370_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call119_367,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv122_371,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_383_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_383_inst_req_0;
      type_cast_383_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_383_inst_req_1;
      type_cast_383_inst_ack_1<= rack(0);
      type_cast_383_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_383_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call124_380,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_384,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_395_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_395_inst_req_0;
      type_cast_395_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_395_inst_req_1;
      type_cast_395_inst_ack_1<= rack(0);
      type_cast_395_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_395_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call128_392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_396,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_408_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_408_inst_req_0;
      type_cast_408_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_408_inst_req_1;
      type_cast_408_inst_ack_1<= rack(0);
      type_cast_408_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_408_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_405,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_409,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_44_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_44_inst_req_0;
      type_cast_44_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_44_inst_req_1;
      type_cast_44_inst_ack_1<= rack(0);
      type_cast_44_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_44_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_41,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_45,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_457_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_457_inst_req_0;
      type_cast_457_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_457_inst_req_1;
      type_cast_457_inst_ack_1<= rack(0);
      type_cast_457_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_457_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp562x_xop_454,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_26_458,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_480_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_480_inst_req_0;
      type_cast_480_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_480_inst_req_1;
      type_cast_480_inst_ack_1<= rack(0);
      type_cast_480_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_480_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext556_631,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_480_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_494_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_494_inst_req_0;
      type_cast_494_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_494_inst_req_1;
      type_cast_494_inst_ack_1<= rack(0);
      type_cast_494_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_494_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call143_491,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv144_495,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_507_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_507_inst_req_0;
      type_cast_507_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_507_inst_req_1;
      type_cast_507_inst_ack_1<= rack(0);
      type_cast_507_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_507_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call147_504,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv149_508,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_525_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_525_inst_req_0;
      type_cast_525_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_525_inst_req_1;
      type_cast_525_inst_ack_1<= rack(0);
      type_cast_525_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_525_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call153_522,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv155_526,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_543_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_543_inst_req_0;
      type_cast_543_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_543_inst_req_1;
      type_cast_543_inst_ack_1<= rack(0);
      type_cast_543_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_543_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call159_540,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv161_544,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_561_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_561_inst_req_0;
      type_cast_561_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_561_inst_req_1;
      type_cast_561_inst_ack_1<= rack(0);
      type_cast_561_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_561_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call165_558,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv167_562,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_579_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_579_inst_req_0;
      type_cast_579_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_579_inst_req_1;
      type_cast_579_inst_ack_1<= rack(0);
      type_cast_579_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_579_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call171_576,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv173_580,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_57_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_57_inst_req_0;
      type_cast_57_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_57_inst_req_1;
      type_cast_57_inst_ack_1<= rack(0);
      type_cast_57_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_57_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_54,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_58,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_597_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_597_inst_req_0;
      type_cast_597_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_597_inst_req_1;
      type_cast_597_inst_ack_1<= rack(0);
      type_cast_597_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_597_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call177_594,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv179_598,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_615_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_615_inst_req_0;
      type_cast_615_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_615_inst_req_1;
      type_cast_615_inst_ack_1<= rack(0);
      type_cast_615_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_615_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call183_612,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv185_616,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_664_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_664_inst_req_0;
      type_cast_664_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_664_inst_req_1;
      type_cast_664_inst_ack_1<= rack(0);
      type_cast_664_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_664_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp548x_xop_661,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_39_665,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_687_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_687_inst_req_0;
      type_cast_687_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_687_inst_req_1;
      type_cast_687_inst_ack_1<= rack(0);
      type_cast_687_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_687_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext540_838,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_687_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_69_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_69_inst_req_0;
      type_cast_69_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_69_inst_req_1;
      type_cast_69_inst_ack_1<= rack(0);
      type_cast_69_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_69_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_66,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_70,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_701_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_701_inst_req_0;
      type_cast_701_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_701_inst_req_1;
      type_cast_701_inst_ack_1<= rack(0);
      type_cast_701_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_701_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call199_698,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_702,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_714_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_714_inst_req_0;
      type_cast_714_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_714_inst_req_1;
      type_cast_714_inst_ack_1<= rack(0);
      type_cast_714_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_714_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call203_711,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv205_715,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_732_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_732_inst_req_0;
      type_cast_732_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_732_inst_req_1;
      type_cast_732_inst_ack_1<= rack(0);
      type_cast_732_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_732_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call209_729,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv211_733,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_750_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_750_inst_req_0;
      type_cast_750_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_750_inst_req_1;
      type_cast_750_inst_ack_1<= rack(0);
      type_cast_750_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_750_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call215_747,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv217_751,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_768_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_768_inst_req_0;
      type_cast_768_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_768_inst_req_1;
      type_cast_768_inst_ack_1<= rack(0);
      type_cast_768_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_768_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call221_765,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv223_769,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_786_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_786_inst_req_0;
      type_cast_786_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_786_inst_req_1;
      type_cast_786_inst_ack_1<= rack(0);
      type_cast_786_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_786_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call227_783,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv229_787,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_804_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_804_inst_req_0;
      type_cast_804_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_804_inst_req_1;
      type_cast_804_inst_ack_1<= rack(0);
      type_cast_804_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_804_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call233_801,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv235_805,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_822_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_822_inst_req_0;
      type_cast_822_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_822_inst_req_1;
      type_cast_822_inst_ack_1<= rack(0);
      type_cast_822_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_822_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call239_819,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv241_823,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_82_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_82_inst_req_0;
      type_cast_82_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_82_inst_req_1;
      type_cast_82_inst_ack_1<= rack(0);
      type_cast_82_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_82_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_79,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_83,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_855_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_855_inst_req_0;
      type_cast_855_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_855_inst_req_1;
      type_cast_855_inst_ack_1<= rack(0);
      type_cast_855_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_855_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add117_364,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv253_856,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_859_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_859_inst_req_0;
      type_cast_859_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_859_inst_req_1;
      type_cast_859_inst_ack_1<= rack(0);
      type_cast_859_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_859_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add126_389,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv255_860,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_863_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_863_inst_req_0;
      type_cast_863_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_863_inst_req_1;
      type_cast_863_inst_ack_1<= rack(0);
      type_cast_863_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_863_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add135_414,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv258_864,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_908_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_908_inst_req_0;
      type_cast_908_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_908_inst_req_1;
      type_cast_908_inst_ack_1<= rack(0);
      type_cast_908_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_908_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp532x_xop_905,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_53_909,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_928_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_928_inst_req_0;
      type_cast_928_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_928_inst_req_1;
      type_cast_928_inst_ack_1<= rack(0);
      type_cast_928_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_928_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext526_950,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_928_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_94_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_94_inst_req_0;
      type_cast_94_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_94_inst_req_1;
      type_cast_94_inst_ack_1<= rack(0);
      type_cast_94_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_94_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_91,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_95,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_972_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_972_inst_req_0;
      type_cast_972_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_972_inst_req_1;
      type_cast_972_inst_ack_1<= rack(0);
      type_cast_972_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_972_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_971_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv276_973,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1368_index_1_rename
    process(R_indvar_1367_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1367_resized;
      ov(13 downto 0) := iv;
      R_indvar_1367_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1368_index_1_resize
    process(indvar_1356) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1356;
      ov := iv(13 downto 0);
      R_indvar_1367_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1368_root_address_inst
    process(array_obj_ref_1368_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1368_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1368_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_486_index_1_rename
    process(R_indvar555_485_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar555_485_resized;
      ov(13 downto 0) := iv;
      R_indvar555_485_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_486_index_1_resize
    process(indvar555_474) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar555_474;
      ov := iv(13 downto 0);
      R_indvar555_485_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_486_root_address_inst
    process(array_obj_ref_486_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_486_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_486_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_693_index_1_rename
    process(R_indvar539_692_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar539_692_resized;
      ov(10 downto 0) := iv;
      R_indvar539_692_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_693_index_1_resize
    process(indvar539_681) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar539_681;
      ov := iv(10 downto 0);
      R_indvar539_692_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_693_root_address_inst
    process(array_obj_ref_693_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_693_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_693_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_937_index_1_rename
    process(R_indvar525_936_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar525_936_resized;
      ov(13 downto 0) := iv;
      R_indvar525_936_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_937_index_1_resize
    process(indvar525_925) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar525_925;
      ov := iv(13 downto 0);
      R_indvar525_936_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_937_root_address_inst
    process(array_obj_ref_937_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_937_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_937_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1373_addr_0
    process(ptr_deref_1373_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1373_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1373_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1373_base_resize
    process(arrayidx432_1370) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx432_1370;
      ov := iv(13 downto 0);
      ptr_deref_1373_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1373_gather_scatter
    process(ptr_deref_1373_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1373_data_0;
      ov(63 downto 0) := iv;
      tmp433_1374 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1373_root_address_inst
    process(ptr_deref_1373_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1373_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1373_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_623_addr_0
    process(ptr_deref_623_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_623_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_623_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_623_base_resize
    process(arrayidx_488) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_488;
      ov := iv(13 downto 0);
      ptr_deref_623_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_623_gather_scatter
    process(add186_621) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add186_621;
      ov(63 downto 0) := iv;
      ptr_deref_623_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_623_root_address_inst
    process(ptr_deref_623_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_623_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_623_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_830_addr_0
    process(ptr_deref_830_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_830_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_830_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_830_base_resize
    process(arrayidx246_695) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx246_695;
      ov := iv(10 downto 0);
      ptr_deref_830_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_830_gather_scatter
    process(add242_828) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add242_828;
      ov(63 downto 0) := iv;
      ptr_deref_830_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_830_root_address_inst
    process(ptr_deref_830_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_830_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_830_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_941_addr_0
    process(ptr_deref_941_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_941_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_941_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_941_base_resize
    process(arrayidx269_939) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx269_939;
      ov := iv(13 downto 0);
      ptr_deref_941_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_941_gather_scatter
    process(type_cast_943_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_943_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_941_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_941_root_address_inst
    process(ptr_deref_941_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_941_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_941_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1312_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264505_880;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1312_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1312_branch_req_0,
          ack0 => if_stmt_1312_branch_ack_0,
          ack1 => if_stmt_1312_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1484_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1483;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1484_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1484_branch_req_0,
          ack0 => if_stmt_1484_branch_ack_0,
          ack1 => if_stmt_1484_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_421_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp513_420;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_421_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_421_branch_req_0,
          ack0 => if_stmt_421_branch_ack_0,
          ack1 => if_stmt_421_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_436_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp194509_435;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_436_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_436_branch_req_0,
          ack0 => if_stmt_436_branch_ack_0,
          ack1 => if_stmt_436_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_637_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_636;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_637_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_637_branch_req_0,
          ack0 => if_stmt_637_branch_ack_0,
          ack1 => if_stmt_637_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_844_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_843;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_844_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_844_branch_req_0,
          ack0 => if_stmt_844_branch_ack_0,
          ack1 => if_stmt_844_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_881_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264505_880;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_881_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_881_branch_req_0,
          ack0 => if_stmt_881_branch_ack_0,
          ack1 => if_stmt_881_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_956_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_955;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_956_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_956_branch_req_0,
          ack0 => if_stmt_956_branch_ack_0,
          ack1 => if_stmt_956_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1335_inst
    process(tmp520_1324) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp520_1324, type_cast_1334_wire_constant, tmp_var);
      tmp520x_xop_1336 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_257_inst
    process(add74_253, shr_241) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add74_253, shr_241, tmp_var);
      add79_258 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_453_inst
    process(shr_241) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr_241, type_cast_452_wire_constant, tmp_var);
      tmp562x_xop_454 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_660_inst
    process(tmp548_649) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp548_649, type_cast_659_wire_constant, tmp_var);
      tmp548x_xop_661 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_904_inst
    process(tmp532_893) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp532_893, type_cast_903_wire_constant, tmp_var);
      tmp532x_xop_905 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1345_inst
    process(iNsTr_196_1340) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_196_1340, type_cast_1344_wire_constant, tmp_var);
      xx_xop_1346 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1477_inst
    process(indvar_1356) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1356, type_cast_1476_wire_constant, tmp_var);
      indvarx_xnext_1478 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_463_inst
    process(iNsTr_26_458) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_26_458, type_cast_462_wire_constant, tmp_var);
      xx_xop571_464 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_630_inst
    process(indvar555_474) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar555_474, type_cast_629_wire_constant, tmp_var);
      indvarx_xnext556_631 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_670_inst
    process(iNsTr_39_665) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_39_665, type_cast_669_wire_constant, tmp_var);
      xx_xop570_671 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_837_inst
    process(indvar539_681) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar539_681, type_cast_836_wire_constant, tmp_var);
      indvarx_xnext540_838 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_914_inst
    process(iNsTr_53_909) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_53_909, type_cast_913_wire_constant, tmp_var);
      xx_xop569_915 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_949_inst
    process(indvar525_925) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar525_925, type_cast_948_wire_constant, tmp_var);
      indvarx_xnext526_950 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_252_inst
    process(iNsTr_14_247) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_14_247, type_cast_251_wire_constant, tmp_var);
      add74_253 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1482_inst
    process(indvarx_xnext_1478, tmp524_1353) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1478, tmp524_1353, tmp_var);
      exitcond1_1483 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_635_inst
    process(indvarx_xnext556_631, tmp567_471) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext556_631, tmp567_471, tmp_var);
      exitcond3_636 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_842_inst
    process(indvarx_xnext540_838, tmp553_678) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext540_838, tmp553_678, tmp_var);
      exitcond2_843 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_954_inst
    process(indvarx_xnext526_950, tmp537_922) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext526_950, tmp537_922, tmp_var);
      exitcond_955 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1050_inst
    process(mul66_235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_235, type_cast_1049_wire_constant, tmp_var);
      shr304_1051 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1106_inst
    process(mul66_235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_235, type_cast_1105_wire_constant, tmp_var);
      shr321_1107 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1162_inst
    process(add79_258) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_258, type_cast_1161_wire_constant, tmp_var);
      shr338_1163 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1323_inst
    process(mul259_874) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_874, type_cast_1322_wire_constant, tmp_var);
      tmp520_1324 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_240_inst
    process(mul66_235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_235, type_cast_239_wire_constant, tmp_var);
      shr_241 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_246_inst
    process(mul66_235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_235, type_cast_245_wire_constant, tmp_var);
      iNsTr_14_247 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_648_inst
    process(mul91_289) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul91_289, type_cast_647_wire_constant, tmp_var);
      tmp548_649 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_892_inst
    process(mul259_874) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_874, type_cast_891_wire_constant, tmp_var);
      tmp532_893 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1221_inst
    process(sub_1212) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1212, type_cast_1220_wire_constant, tmp_var);
      shr364_1222 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1231_inst
    process(sub_1212) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1212, type_cast_1230_wire_constant, tmp_var);
      shr370_1232 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1241_inst
    process(sub_1212) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1212, type_cast_1240_wire_constant, tmp_var);
      shr376_1242 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1251_inst
    process(sub_1212) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1212, type_cast_1250_wire_constant, tmp_var);
      shr382_1252 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1261_inst
    process(sub_1212) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1212, type_cast_1260_wire_constant, tmp_var);
      shr388_1262 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1271_inst
    process(sub_1212) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1212, type_cast_1270_wire_constant, tmp_var);
      shr394_1272 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1281_inst
    process(sub_1212) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1212, type_cast_1280_wire_constant, tmp_var);
      shr400_1282 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1383_inst
    process(tmp433_1374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1374, type_cast_1382_wire_constant, tmp_var);
      shr440_1384 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1393_inst
    process(tmp433_1374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1374, type_cast_1392_wire_constant, tmp_var);
      shr446_1394 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1403_inst
    process(tmp433_1374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1374, type_cast_1402_wire_constant, tmp_var);
      shr452_1404 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1413_inst
    process(tmp433_1374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1374, type_cast_1412_wire_constant, tmp_var);
      shr458_1414 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1423_inst
    process(tmp433_1374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1374, type_cast_1422_wire_constant, tmp_var);
      shr464_1424 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1433_inst
    process(tmp433_1374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1374, type_cast_1432_wire_constant, tmp_var);
      shr470_1434 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1443_inst
    process(tmp433_1374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1374, type_cast_1442_wire_constant, tmp_var);
      shr476_1444 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_229_inst
    process(conv63_221, conv61_217) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv63_221, conv61_217, tmp_var);
      mul_230 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_234_inst
    process(mul_230, conv65_225) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_230, conv65_225, tmp_var);
      mul66_235 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_278_inst
    process(conv84_266, conv82_262) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv84_266, conv82_262, tmp_var);
      mul85_279 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_283_inst
    process(mul85_279, conv87_270) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul85_279, conv87_270, tmp_var);
      mul88_284 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_288_inst
    process(mul88_284, conv90_274) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul88_284, conv90_274, tmp_var);
      mul91_289 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_868_inst
    process(conv255_860, conv253_856) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv255_860, conv253_856, tmp_var);
      mul256_869 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_873_inst
    process(mul256_869, conv258_864) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul256_869, conv258_864, tmp_var);
      mul259_874 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_112_inst
    process(shl18_101, conv20_108) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_101, conv20_108, tmp_var);
      add21_113 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_137_inst
    process(shl27_126, conv29_133) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_126, conv29_133, tmp_var);
      add30_138 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_162_inst
    process(shl36_151, conv38_158) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_151, conv38_158, tmp_var);
      add39_163 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_187_inst
    process(shl45_176, conv47_183) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_176, conv47_183, tmp_var);
      add48_188 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_212_inst
    process(shl54_201, conv56_208) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_201, conv56_208, tmp_var);
      add57_213 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_313_inst
    process(shl96_302, conv98_309) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl96_302, conv98_309, tmp_var);
      add99_314 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_338_inst
    process(shl105_327, conv107_334) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl105_327, conv107_334, tmp_var);
      add108_339 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_363_inst
    process(shl114_352, conv116_359) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl114_352, conv116_359, tmp_var);
      add117_364 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_388_inst
    process(shl123_377, conv125_384) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl123_377, conv125_384, tmp_var);
      add126_389 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_413_inst
    process(shl132_402, conv134_409) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_402, conv134_409, tmp_var);
      add135_414 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_62_inst
    process(shl_51, conv3_58) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_51, conv3_58, tmp_var);
      add_63 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_87_inst
    process(shl9_76, conv11_83) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_76, conv11_83, tmp_var);
      add12_88 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_512_inst
    process(shl146_501, conv149_508) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl146_501, conv149_508, tmp_var);
      add150_513 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_530_inst
    process(shl152_519, conv155_526) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl152_519, conv155_526, tmp_var);
      add156_531 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_548_inst
    process(shl158_537, conv161_544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl158_537, conv161_544, tmp_var);
      add162_549 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_566_inst
    process(shl164_555, conv167_562) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl164_555, conv167_562, tmp_var);
      add168_567 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_584_inst
    process(shl170_573, conv173_580) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl170_573, conv173_580, tmp_var);
      add174_585 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_602_inst
    process(shl176_591, conv179_598) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl176_591, conv179_598, tmp_var);
      add180_603 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_620_inst
    process(shl182_609, conv185_616) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl182_609, conv185_616, tmp_var);
      add186_621 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_719_inst
    process(shl202_708, conv205_715) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl202_708, conv205_715, tmp_var);
      add206_720 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_737_inst
    process(shl208_726, conv211_733) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl208_726, conv211_733, tmp_var);
      add212_738 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_755_inst
    process(shl214_744, conv217_751) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl214_744, conv217_751, tmp_var);
      add218_756 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_773_inst
    process(shl220_762, conv223_769) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl220_762, conv223_769, tmp_var);
      add224_774 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_791_inst
    process(shl226_780, conv229_787) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl226_780, conv229_787, tmp_var);
      add230_792 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_809_inst
    process(shl232_798, conv235_805) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl232_798, conv235_805, tmp_var);
      add236_810 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_827_inst
    process(shl238_816, conv241_823) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl238_816, conv241_823, tmp_var);
      add242_828 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_100_inst
    process(conv17_95) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_95, type_cast_99_wire_constant, tmp_var);
      shl18_101 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_125_inst
    process(conv26_120) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_120, type_cast_124_wire_constant, tmp_var);
      shl27_126 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_150_inst
    process(conv35_145) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_145, type_cast_149_wire_constant, tmp_var);
      shl36_151 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_175_inst
    process(conv44_170) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_170, type_cast_174_wire_constant, tmp_var);
      shl45_176 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_200_inst
    process(conv53_195) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_195, type_cast_199_wire_constant, tmp_var);
      shl54_201 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_301_inst
    process(conv95_296) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv95_296, type_cast_300_wire_constant, tmp_var);
      shl96_302 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_326_inst
    process(conv104_321) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv104_321, type_cast_325_wire_constant, tmp_var);
      shl105_327 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_351_inst
    process(conv113_346) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv113_346, type_cast_350_wire_constant, tmp_var);
      shl114_352 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_376_inst
    process(conv122_371) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv122_371, type_cast_375_wire_constant, tmp_var);
      shl123_377 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_401_inst
    process(conv131_396) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv131_396, type_cast_400_wire_constant, tmp_var);
      shl132_402 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_50_inst
    process(conv1_45) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_45, type_cast_49_wire_constant, tmp_var);
      shl_51 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_75_inst
    process(conv8_70) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_70, type_cast_74_wire_constant, tmp_var);
      shl9_76 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_500_inst
    process(conv144_495) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv144_495, type_cast_499_wire_constant, tmp_var);
      shl146_501 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_518_inst
    process(add150_513) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add150_513, type_cast_517_wire_constant, tmp_var);
      shl152_519 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_536_inst
    process(add156_531) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add156_531, type_cast_535_wire_constant, tmp_var);
      shl158_537 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_554_inst
    process(add162_549) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add162_549, type_cast_553_wire_constant, tmp_var);
      shl164_555 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_572_inst
    process(add168_567) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add168_567, type_cast_571_wire_constant, tmp_var);
      shl170_573 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_590_inst
    process(add174_585) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add174_585, type_cast_589_wire_constant, tmp_var);
      shl176_591 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_608_inst
    process(add180_603) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add180_603, type_cast_607_wire_constant, tmp_var);
      shl182_609 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_707_inst
    process(conv200_702) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv200_702, type_cast_706_wire_constant, tmp_var);
      shl202_708 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_725_inst
    process(add206_720) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add206_720, type_cast_724_wire_constant, tmp_var);
      shl208_726 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_743_inst
    process(add212_738) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add212_738, type_cast_742_wire_constant, tmp_var);
      shl214_744 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_761_inst
    process(add218_756) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add218_756, type_cast_760_wire_constant, tmp_var);
      shl220_762 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_779_inst
    process(add224_774) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add224_774, type_cast_778_wire_constant, tmp_var);
      shl226_780 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_797_inst
    process(add230_792) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add230_792, type_cast_796_wire_constant, tmp_var);
      shl232_798 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_815_inst
    process(add236_810) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add236_810, type_cast_814_wire_constant, tmp_var);
      shl238_816 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1211_inst
    process(conv355_1207, conv276_973) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv355_1207, conv276_973, tmp_var);
      sub_1212 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1329_inst
    process(tmp520_1324) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp520_1324, type_cast_1328_wire_constant, tmp_var);
      tmp521_1330 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_419_inst
    process(mul66_235) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul66_235, type_cast_418_wire_constant, tmp_var);
      cmp513_420 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_434_inst
    process(mul91_289) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul91_289, type_cast_433_wire_constant, tmp_var);
      cmp194509_435 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_447_inst
    process(shr_241) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_241, type_cast_446_wire_constant, tmp_var);
      tmp563_448 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_654_inst
    process(tmp548_649) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp548_649, type_cast_653_wire_constant, tmp_var);
      tmp549_655 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_879_inst
    process(mul259_874) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul259_874, type_cast_878_wire_constant, tmp_var);
      cmp264505_880 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_898_inst
    process(tmp532_893) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp532_893, type_cast_897_wire_constant, tmp_var);
      tmp533_899 <= tmp_var; --
    end process;
    -- shared split operator group (107) : array_obj_ref_1368_index_offset 
    ApIntAdd_group_107: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1367_scaled;
      array_obj_ref_1368_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1368_index_offset_req_0;
      array_obj_ref_1368_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1368_index_offset_req_1;
      array_obj_ref_1368_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_107_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_107_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_107",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 107
    -- shared split operator group (108) : array_obj_ref_486_index_offset 
    ApIntAdd_group_108: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar555_485_scaled;
      array_obj_ref_486_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_486_index_offset_req_0;
      array_obj_ref_486_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_486_index_offset_req_1;
      array_obj_ref_486_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_108_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_108_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_108",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 108
    -- shared split operator group (109) : array_obj_ref_693_index_offset 
    ApIntAdd_group_109: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar539_692_scaled;
      array_obj_ref_693_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_693_index_offset_req_0;
      array_obj_ref_693_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_693_index_offset_req_1;
      array_obj_ref_693_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_109_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_109_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_109",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100010",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 109
    -- shared split operator group (110) : array_obj_ref_937_index_offset 
    ApIntAdd_group_110: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar525_936_scaled;
      array_obj_ref_937_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_937_index_offset_req_0;
      array_obj_ref_937_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_937_index_offset_req_1;
      array_obj_ref_937_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_110_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_110_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_110",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 110
    -- unary operator type_cast_1205_inst
    process(call354_1202) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call354_1202, tmp_var);
      type_cast_1205_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_971_inst
    process(call275_967) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call275_967, tmp_var);
      type_cast_971_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1373_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1373_load_0_req_0;
      ptr_deref_1373_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1373_load_0_req_1;
      ptr_deref_1373_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1373_word_address_0;
      ptr_deref_1373_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(13 downto 0),
          mtag => memory_space_2_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_623_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_623_store_0_req_0;
      ptr_deref_623_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_623_store_0_req_1;
      ptr_deref_623_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_623_word_address_0;
      data_in <= ptr_deref_623_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_830_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_830_store_0_req_0;
      ptr_deref_830_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_830_store_0_req_1;
      ptr_deref_830_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_830_word_address_0;
      data_in <= ptr_deref_830_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(10 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_941_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_941_store_0_req_0;
      ptr_deref_941_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_941_store_0_req_1;
      ptr_deref_941_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_941_word_address_0;
      data_in <= ptr_deref_941_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_Block0_done_1189_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1189_inst_req_0;
      RPIPE_Block0_done_1189_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1189_inst_req_1;
      RPIPE_Block0_done_1189_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call346_1190 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1192_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1192_inst_req_0;
      RPIPE_Block1_done_1192_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1192_inst_req_1;
      RPIPE_Block1_done_1192_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call348_1193 <= data_out(15 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1195_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1195_inst_req_0;
      RPIPE_Block2_done_1195_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1195_inst_req_1;
      RPIPE_Block2_done_1195_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call350_1196 <= data_out(15 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1198_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1198_inst_req_0;
      RPIPE_Block3_done_1198_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1198_inst_req_1;
      RPIPE_Block3_done_1198_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call352_1199 <= data_out(15 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_ConvTranspose_input_pipe_53_inst RPIPE_ConvTranspose_input_pipe_40_inst RPIPE_ConvTranspose_input_pipe_710_inst RPIPE_ConvTranspose_input_pipe_128_inst RPIPE_ConvTranspose_input_pipe_697_inst RPIPE_ConvTranspose_input_pipe_818_inst RPIPE_ConvTranspose_input_pipe_782_inst RPIPE_ConvTranspose_input_pipe_728_inst RPIPE_ConvTranspose_input_pipe_153_inst RPIPE_ConvTranspose_input_pipe_178_inst RPIPE_ConvTranspose_input_pipe_140_inst RPIPE_ConvTranspose_input_pipe_800_inst RPIPE_ConvTranspose_input_pipe_115_inst RPIPE_ConvTranspose_input_pipe_78_inst RPIPE_ConvTranspose_input_pipe_746_inst RPIPE_ConvTranspose_input_pipe_165_inst RPIPE_ConvTranspose_input_pipe_764_inst RPIPE_ConvTranspose_input_pipe_90_inst RPIPE_ConvTranspose_input_pipe_103_inst RPIPE_ConvTranspose_input_pipe_65_inst RPIPE_ConvTranspose_input_pipe_190_inst RPIPE_ConvTranspose_input_pipe_203_inst RPIPE_ConvTranspose_input_pipe_291_inst RPIPE_ConvTranspose_input_pipe_304_inst RPIPE_ConvTranspose_input_pipe_316_inst RPIPE_ConvTranspose_input_pipe_329_inst RPIPE_ConvTranspose_input_pipe_341_inst RPIPE_ConvTranspose_input_pipe_354_inst RPIPE_ConvTranspose_input_pipe_366_inst RPIPE_ConvTranspose_input_pipe_379_inst RPIPE_ConvTranspose_input_pipe_391_inst RPIPE_ConvTranspose_input_pipe_404_inst RPIPE_ConvTranspose_input_pipe_490_inst RPIPE_ConvTranspose_input_pipe_503_inst RPIPE_ConvTranspose_input_pipe_521_inst RPIPE_ConvTranspose_input_pipe_539_inst RPIPE_ConvTranspose_input_pipe_557_inst RPIPE_ConvTranspose_input_pipe_575_inst RPIPE_ConvTranspose_input_pipe_593_inst RPIPE_ConvTranspose_input_pipe_611_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(319 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 39 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 39 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 39 downto 0);
      signal guard_vector : std_logic_vector( 39 downto 0);
      constant outBUFs : IntegerArray(39 downto 0) := (39 => 1, 38 => 1, 37 => 1, 36 => 1, 35 => 1, 34 => 1, 33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(39 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false, 35 => false, 36 => false, 37 => false, 38 => false, 39 => false);
      constant guardBuffering: IntegerArray(39 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2, 35 => 2, 36 => 2, 37 => 2, 38 => 2, 39 => 2);
      -- 
    begin -- 
      reqL_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_53_inst_req_0;
      reqL_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_40_inst_req_0;
      reqL_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_710_inst_req_0;
      reqL_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_128_inst_req_0;
      reqL_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_697_inst_req_0;
      reqL_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_818_inst_req_0;
      reqL_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_782_inst_req_0;
      reqL_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_728_inst_req_0;
      reqL_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_153_inst_req_0;
      reqL_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_178_inst_req_0;
      reqL_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_140_inst_req_0;
      reqL_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_800_inst_req_0;
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_115_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_78_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_746_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_165_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_764_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_90_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_103_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_65_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_190_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_203_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_291_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_304_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_316_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_329_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_341_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_354_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_366_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_379_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_391_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_404_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_490_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_503_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_521_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_539_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_557_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_575_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_593_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_611_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_53_inst_ack_0 <= ackL_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_40_inst_ack_0 <= ackL_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_710_inst_ack_0 <= ackL_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_128_inst_ack_0 <= ackL_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_697_inst_ack_0 <= ackL_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_818_inst_ack_0 <= ackL_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_782_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_728_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_153_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_178_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_140_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_800_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_115_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_78_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_746_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_165_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_764_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_90_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_103_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_65_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_190_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_203_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_291_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_304_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_316_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_329_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_341_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_354_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_366_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_379_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_391_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_404_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_490_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_503_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_521_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_539_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_557_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_575_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_593_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_611_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_53_inst_req_1;
      reqR_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_40_inst_req_1;
      reqR_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_710_inst_req_1;
      reqR_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_128_inst_req_1;
      reqR_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_697_inst_req_1;
      reqR_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_818_inst_req_1;
      reqR_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_782_inst_req_1;
      reqR_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_728_inst_req_1;
      reqR_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_153_inst_req_1;
      reqR_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_178_inst_req_1;
      reqR_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_140_inst_req_1;
      reqR_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_800_inst_req_1;
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_115_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_78_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_746_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_165_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_764_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_90_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_103_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_65_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_190_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_203_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_291_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_304_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_316_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_329_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_341_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_354_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_366_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_379_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_391_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_404_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_490_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_503_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_521_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_539_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_557_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_575_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_593_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_611_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_53_inst_ack_1 <= ackR_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_40_inst_ack_1 <= ackR_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_710_inst_ack_1 <= ackR_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_128_inst_ack_1 <= ackR_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_697_inst_ack_1 <= ackR_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_818_inst_ack_1 <= ackR_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_782_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_728_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_153_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_178_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_140_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_800_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_115_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_78_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_746_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_165_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_764_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_90_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_103_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_65_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_190_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_203_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_291_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_304_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_316_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_329_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_341_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_354_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_366_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_379_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_391_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_404_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_490_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_503_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_521_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_539_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_557_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_575_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_593_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_611_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      call2_54 <= data_out(319 downto 312);
      call_41 <= data_out(311 downto 304);
      call203_711 <= data_out(303 downto 296);
      call28_129 <= data_out(295 downto 288);
      call199_698 <= data_out(287 downto 280);
      call239_819 <= data_out(279 downto 272);
      call227_783 <= data_out(271 downto 264);
      call209_729 <= data_out(263 downto 256);
      call37_154 <= data_out(255 downto 248);
      call46_179 <= data_out(247 downto 240);
      call32_141 <= data_out(239 downto 232);
      call233_801 <= data_out(231 downto 224);
      call23_116 <= data_out(223 downto 216);
      call10_79 <= data_out(215 downto 208);
      call215_747 <= data_out(207 downto 200);
      call41_166 <= data_out(199 downto 192);
      call221_765 <= data_out(191 downto 184);
      call14_91 <= data_out(183 downto 176);
      call19_104 <= data_out(175 downto 168);
      call5_66 <= data_out(167 downto 160);
      call50_191 <= data_out(159 downto 152);
      call55_204 <= data_out(151 downto 144);
      call92_292 <= data_out(143 downto 136);
      call97_305 <= data_out(135 downto 128);
      call101_317 <= data_out(127 downto 120);
      call106_330 <= data_out(119 downto 112);
      call110_342 <= data_out(111 downto 104);
      call115_355 <= data_out(103 downto 96);
      call119_367 <= data_out(95 downto 88);
      call124_380 <= data_out(87 downto 80);
      call128_392 <= data_out(79 downto 72);
      call133_405 <= data_out(71 downto 64);
      call143_491 <= data_out(63 downto 56);
      call147_504 <= data_out(55 downto 48);
      call153_522 <= data_out(47 downto 40);
      call159_540 <= data_out(39 downto 32);
      call165_558 <= data_out(31 downto 24);
      call171_576 <= data_out(23 downto 16);
      call177_594 <= data_out(15 downto 8);
      call183_612 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_4_gI", nreqs => 40, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_4: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_4", data_width => 8,  num_reqs => 40,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared outport operator group (0) : WPIPE_Block0_start_1013_inst WPIPE_Block0_start_975_inst WPIPE_Block0_start_978_inst WPIPE_Block0_start_981_inst WPIPE_Block0_start_990_inst WPIPE_Block0_start_993_inst WPIPE_Block0_start_996_inst WPIPE_Block0_start_999_inst WPIPE_Block0_start_984_inst WPIPE_Block0_start_1002_inst WPIPE_Block0_start_987_inst WPIPE_Block0_start_1006_inst WPIPE_Block0_start_1010_inst WPIPE_Block0_start_1016_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block0_start_1013_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block0_start_975_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block0_start_978_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block0_start_981_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block0_start_990_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block0_start_993_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block0_start_996_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block0_start_999_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block0_start_984_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block0_start_1002_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block0_start_987_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block0_start_1006_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block0_start_1010_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block0_start_1016_inst_req_0;
      WPIPE_Block0_start_1013_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block0_start_975_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block0_start_978_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block0_start_981_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block0_start_990_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block0_start_993_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block0_start_996_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block0_start_999_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block0_start_984_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block0_start_1002_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block0_start_987_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block0_start_1006_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block0_start_1010_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block0_start_1016_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block0_start_1013_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block0_start_975_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block0_start_978_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block0_start_981_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block0_start_990_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block0_start_993_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block0_start_996_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block0_start_999_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block0_start_984_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block0_start_1002_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block0_start_987_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block0_start_1006_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block0_start_1010_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block0_start_1016_inst_req_1;
      WPIPE_Block0_start_1013_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block0_start_975_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block0_start_978_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block0_start_981_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block0_start_990_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block0_start_993_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block0_start_996_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block0_start_999_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block0_start_984_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block0_start_1002_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block0_start_987_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block0_start_1006_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block0_start_1010_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block0_start_1016_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add126_389 & add_63 & add12_88 & add21_113 & add48_188 & add57_213 & add99_314 & add108_339 & add30_138 & type_cast_1004_wire_constant & add39_163 & type_cast_1008_wire_constant & add117_364 & add135_414;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_1056_inst WPIPE_Block1_start_1022_inst WPIPE_Block1_start_1063_inst WPIPE_Block1_start_1066_inst WPIPE_Block1_start_1031_inst WPIPE_Block1_start_1034_inst WPIPE_Block1_start_1069_inst WPIPE_Block1_start_1025_inst WPIPE_Block1_start_1072_inst WPIPE_Block1_start_1037_inst WPIPE_Block1_start_1019_inst WPIPE_Block1_start_1028_inst WPIPE_Block1_start_1040_inst WPIPE_Block1_start_1043_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block1_start_1056_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block1_start_1022_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block1_start_1063_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block1_start_1066_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block1_start_1031_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block1_start_1034_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block1_start_1069_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block1_start_1025_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block1_start_1072_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block1_start_1037_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block1_start_1019_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block1_start_1028_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block1_start_1040_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block1_start_1043_inst_req_0;
      WPIPE_Block1_start_1056_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block1_start_1022_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block1_start_1063_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block1_start_1066_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block1_start_1031_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block1_start_1034_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block1_start_1069_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block1_start_1025_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block1_start_1072_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block1_start_1037_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block1_start_1019_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block1_start_1028_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block1_start_1040_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block1_start_1043_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block1_start_1056_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block1_start_1022_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block1_start_1063_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block1_start_1066_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block1_start_1031_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block1_start_1034_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block1_start_1069_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block1_start_1025_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block1_start_1072_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block1_start_1037_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block1_start_1019_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block1_start_1028_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block1_start_1040_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block1_start_1043_inst_req_1;
      WPIPE_Block1_start_1056_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block1_start_1022_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block1_start_1063_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block1_start_1066_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block1_start_1031_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block1_start_1034_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block1_start_1069_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block1_start_1025_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block1_start_1072_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block1_start_1037_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block1_start_1019_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block1_start_1028_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block1_start_1040_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block1_start_1043_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= conv305_1055 & add12_88 & conv307_1062 & add117_364 & add39_163 & add48_188 & add126_389 & add21_113 & add135_414 & add57_213 & add_63 & add30_138 & add99_314 & add108_339;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1090_inst WPIPE_Block2_start_1112_inst WPIPE_Block2_start_1128_inst WPIPE_Block2_start_1087_inst WPIPE_Block2_start_1093_inst WPIPE_Block2_start_1096_inst WPIPE_Block2_start_1084_inst WPIPE_Block2_start_1099_inst WPIPE_Block2_start_1075_inst WPIPE_Block2_start_1078_inst WPIPE_Block2_start_1081_inst WPIPE_Block2_start_1119_inst WPIPE_Block2_start_1122_inst WPIPE_Block2_start_1125_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block2_start_1090_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block2_start_1112_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block2_start_1128_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block2_start_1087_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block2_start_1093_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block2_start_1096_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block2_start_1084_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block2_start_1099_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block2_start_1075_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block2_start_1078_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block2_start_1081_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block2_start_1119_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block2_start_1122_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block2_start_1125_inst_req_0;
      WPIPE_Block2_start_1090_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block2_start_1112_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block2_start_1128_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block2_start_1087_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block2_start_1093_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block2_start_1096_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block2_start_1084_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block2_start_1099_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block2_start_1075_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block2_start_1078_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block2_start_1081_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block2_start_1119_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block2_start_1122_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block2_start_1125_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block2_start_1090_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block2_start_1112_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block2_start_1128_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block2_start_1087_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block2_start_1093_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block2_start_1096_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block2_start_1084_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block2_start_1099_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block2_start_1075_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block2_start_1078_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block2_start_1081_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block2_start_1119_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block2_start_1122_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block2_start_1125_inst_req_1;
      WPIPE_Block2_start_1090_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block2_start_1112_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block2_start_1128_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block2_start_1087_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block2_start_1093_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block2_start_1096_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block2_start_1084_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block2_start_1099_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block2_start_1075_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block2_start_1078_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block2_start_1081_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block2_start_1119_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block2_start_1122_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block2_start_1125_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add48_188 & conv322_1111 & add135_414 & add39_163 & add57_213 & add99_314 & add30_138 & add108_339 & add_63 & add12_88 & add21_113 & conv324_1118 & add117_364 & add126_389;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1134_inst WPIPE_Block3_start_1149_inst WPIPE_Block3_start_1178_inst WPIPE_Block3_start_1131_inst WPIPE_Block3_start_1137_inst WPIPE_Block3_start_1143_inst WPIPE_Block3_start_1152_inst WPIPE_Block3_start_1140_inst WPIPE_Block3_start_1168_inst WPIPE_Block3_start_1181_inst WPIPE_Block3_start_1155_inst WPIPE_Block3_start_1146_inst WPIPE_Block3_start_1184_inst WPIPE_Block3_start_1175_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block3_start_1134_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block3_start_1149_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block3_start_1178_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block3_start_1131_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block3_start_1137_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block3_start_1143_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block3_start_1152_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block3_start_1140_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block3_start_1168_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block3_start_1181_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block3_start_1155_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block3_start_1146_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block3_start_1184_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block3_start_1175_inst_req_0;
      WPIPE_Block3_start_1134_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block3_start_1149_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block3_start_1178_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block3_start_1131_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block3_start_1137_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block3_start_1143_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block3_start_1152_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block3_start_1140_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block3_start_1168_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block3_start_1181_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block3_start_1155_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block3_start_1146_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block3_start_1184_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block3_start_1175_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block3_start_1134_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block3_start_1149_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block3_start_1178_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block3_start_1131_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block3_start_1137_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block3_start_1143_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block3_start_1152_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block3_start_1140_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block3_start_1168_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block3_start_1181_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block3_start_1155_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block3_start_1146_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block3_start_1184_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block3_start_1175_inst_req_1;
      WPIPE_Block3_start_1134_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block3_start_1149_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block3_start_1178_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block3_start_1131_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block3_start_1137_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block3_start_1143_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block3_start_1152_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block3_start_1140_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block3_start_1168_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block3_start_1181_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block3_start_1155_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block3_start_1146_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block3_start_1184_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block3_start_1175_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add12_88 & add57_213 & add117_364 & add_63 & add21_113 & add39_163 & add99_314 & add30_138 & conv339_1167 & add126_389 & add108_339 & add48_188 & add135_414 & conv341_1174;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_ConvTranspose_output_pipe_1302_inst WPIPE_ConvTranspose_output_pipe_1299_inst WPIPE_ConvTranspose_output_pipe_1296_inst WPIPE_ConvTranspose_output_pipe_1287_inst WPIPE_ConvTranspose_output_pipe_1293_inst WPIPE_ConvTranspose_output_pipe_1290_inst WPIPE_ConvTranspose_output_pipe_1308_inst WPIPE_ConvTranspose_output_pipe_1305_inst WPIPE_ConvTranspose_output_pipe_1449_inst WPIPE_ConvTranspose_output_pipe_1452_inst WPIPE_ConvTranspose_output_pipe_1455_inst WPIPE_ConvTranspose_output_pipe_1458_inst WPIPE_ConvTranspose_output_pipe_1461_inst WPIPE_ConvTranspose_output_pipe_1464_inst WPIPE_ConvTranspose_output_pipe_1467_inst WPIPE_ConvTranspose_output_pipe_1470_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 15 downto 0);
      signal update_req, update_ack : BooleanArray( 15 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 15 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      sample_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1302_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1299_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1296_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1287_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1293_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1290_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1308_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1305_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1449_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1452_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1455_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1458_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1461_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1464_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1467_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1470_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1302_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1299_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1296_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1287_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1293_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1290_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1308_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1305_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1449_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1452_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1455_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1458_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1461_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1464_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1467_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1470_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1302_inst_req_1;
      update_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1299_inst_req_1;
      update_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1296_inst_req_1;
      update_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1287_inst_req_1;
      update_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1293_inst_req_1;
      update_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1290_inst_req_1;
      update_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1308_inst_req_1;
      update_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1305_inst_req_1;
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1449_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1452_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1455_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1458_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1461_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1464_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1467_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1470_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1302_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1299_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1296_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1287_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1293_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1290_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1308_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1305_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1449_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1452_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1455_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1458_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1461_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1464_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1467_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1470_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      data_in <= conv373_1236 & conv379_1246 & conv385_1256 & conv403_1286 & conv391_1266 & conv397_1276 & conv361_1216 & conv367_1226 & conv479_1448 & conv473_1438 & conv467_1428 & conv461_1418 & conv455_1408 & conv449_1398 & conv443_1388 & conv437_1378;
      ConvTranspose_output_pipe_write_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_4_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_4: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 16, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared call operator group (0) : call_stmt_1202_call call_stmt_967_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1202_call_req_0;
      reqL_unguarded(0) <= call_stmt_967_call_req_0;
      call_stmt_1202_call_ack_0 <= ackL_unguarded(1);
      call_stmt_967_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1202_call_req_1;
      reqR_unguarded(0) <= call_stmt_967_call_req_1;
      call_stmt_1202_call_ack_1 <= ackR_unguarded(1);
      call_stmt_967_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call354_1202 <= data_out(127 downto 64);
      call275_967 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_3763_start: Boolean;
  signal convTransposeA_CP_3763_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1822_inst_req_1 : boolean;
  signal type_cast_1613_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1515_inst_ack_1 : boolean;
  signal type_cast_1822_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1540_inst_req_0 : boolean;
  signal type_cast_1531_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1509_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1552_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1506_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1500_inst_ack_1 : boolean;
  signal phi_stmt_1607_req_1 : boolean;
  signal RPIPE_Block0_start_1506_inst_ack_1 : boolean;
  signal type_cast_1634_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1503_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1500_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1552_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1540_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1555_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1527_inst_req_1 : boolean;
  signal type_cast_1634_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1506_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1527_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1555_inst_req_0 : boolean;
  signal phi_stmt_1607_ack_0 : boolean;
  signal RPIPE_Block0_start_1558_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1524_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1509_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1527_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1524_inst_ack_0 : boolean;
  signal type_cast_1531_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1527_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1503_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1518_inst_req_0 : boolean;
  signal phi_stmt_1823_ack_0 : boolean;
  signal RPIPE_Block0_start_1518_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1540_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1521_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1558_inst_req_1 : boolean;
  signal type_cast_1826_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1503_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1555_inst_ack_0 : boolean;
  signal phi_stmt_1621_req_0 : boolean;
  signal RPIPE_Block0_start_1509_inst_ack_1 : boolean;
  signal type_cast_1531_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1515_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1503_inst_ack_0 : boolean;
  signal phi_stmt_1816_req_0 : boolean;
  signal RPIPE_Block0_start_1515_inst_ack_0 : boolean;
  signal type_cast_1634_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1521_inst_req_1 : boolean;
  signal phi_stmt_1621_ack_0 : boolean;
  signal RPIPE_Block0_start_1518_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1512_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1540_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1521_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1555_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1521_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1512_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1558_inst_req_0 : boolean;
  signal phi_stmt_1823_req_0 : boolean;
  signal RPIPE_Block0_start_1558_inst_ack_0 : boolean;
  signal type_cast_1531_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1515_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1518_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1506_inst_req_1 : boolean;
  signal type_cast_1613_inst_req_1 : boolean;
  signal phi_stmt_1614_ack_0 : boolean;
  signal RPIPE_Block0_start_1552_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1500_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1500_inst_ack_0 : boolean;
  signal phi_stmt_1628_ack_0 : boolean;
  signal phi_stmt_1607_req_0 : boolean;
  signal type_cast_1613_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1512_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1552_inst_req_0 : boolean;
  signal type_cast_1589_inst_ack_1 : boolean;
  signal type_cast_1589_inst_req_1 : boolean;
  signal type_cast_1589_inst_req_0 : boolean;
  signal type_cast_1589_inst_ack_0 : boolean;
  signal type_cast_1634_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1509_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1512_inst_ack_0 : boolean;
  signal type_cast_1585_inst_req_1 : boolean;
  signal type_cast_1826_inst_req_1 : boolean;
  signal type_cast_1585_inst_ack_1 : boolean;
  signal type_cast_1585_inst_ack_0 : boolean;
  signal type_cast_1544_inst_ack_1 : boolean;
  signal phi_stmt_1628_req_1 : boolean;
  signal type_cast_1585_inst_req_0 : boolean;
  signal type_cast_1544_inst_req_1 : boolean;
  signal type_cast_1822_inst_req_0 : boolean;
  signal phi_stmt_1816_ack_0 : boolean;
  signal RPIPE_Block0_start_1524_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1524_inst_req_1 : boolean;
  signal type_cast_1544_inst_ack_0 : boolean;
  signal type_cast_1544_inst_req_0 : boolean;
  signal type_cast_1822_inst_ack_0 : boolean;
  signal type_cast_1593_inst_req_0 : boolean;
  signal type_cast_1826_inst_ack_0 : boolean;
  signal type_cast_1593_inst_ack_0 : boolean;
  signal type_cast_1826_inst_req_0 : boolean;
  signal type_cast_1593_inst_req_1 : boolean;
  signal type_cast_1593_inst_ack_1 : boolean;
  signal type_cast_1597_inst_req_0 : boolean;
  signal type_cast_1597_inst_ack_0 : boolean;
  signal type_cast_1597_inst_req_1 : boolean;
  signal type_cast_1597_inst_ack_1 : boolean;
  signal phi_stmt_1621_req_1 : boolean;
  signal phi_stmt_1823_req_1 : boolean;
  signal type_cast_1669_inst_req_0 : boolean;
  signal type_cast_1669_inst_ack_0 : boolean;
  signal type_cast_1669_inst_req_1 : boolean;
  signal type_cast_1669_inst_ack_1 : boolean;
  signal type_cast_1828_inst_ack_1 : boolean;
  signal type_cast_1828_inst_req_1 : boolean;
  signal type_cast_1627_inst_ack_1 : boolean;
  signal type_cast_1673_inst_req_0 : boolean;
  signal type_cast_1673_inst_ack_0 : boolean;
  signal type_cast_1673_inst_req_1 : boolean;
  signal type_cast_1673_inst_ack_1 : boolean;
  signal type_cast_1627_inst_req_1 : boolean;
  signal type_cast_1828_inst_ack_0 : boolean;
  signal type_cast_1677_inst_req_0 : boolean;
  signal type_cast_1677_inst_ack_0 : boolean;
  signal type_cast_1613_inst_req_0 : boolean;
  signal type_cast_1677_inst_req_1 : boolean;
  signal type_cast_1677_inst_ack_1 : boolean;
  signal type_cast_1828_inst_req_0 : boolean;
  signal type_cast_1707_inst_req_0 : boolean;
  signal type_cast_1707_inst_ack_0 : boolean;
  signal type_cast_1707_inst_req_1 : boolean;
  signal type_cast_1707_inst_ack_1 : boolean;
  signal type_cast_1627_inst_ack_0 : boolean;
  signal type_cast_1627_inst_req_0 : boolean;
  signal array_obj_ref_1713_index_offset_req_0 : boolean;
  signal phi_stmt_1829_req_0 : boolean;
  signal array_obj_ref_1713_index_offset_ack_0 : boolean;
  signal array_obj_ref_1713_index_offset_req_1 : boolean;
  signal type_cast_1832_inst_ack_1 : boolean;
  signal array_obj_ref_1713_index_offset_ack_1 : boolean;
  signal phi_stmt_1816_req_1 : boolean;
  signal type_cast_1832_inst_req_1 : boolean;
  signal phi_stmt_1628_req_0 : boolean;
  signal addr_of_1714_final_reg_req_0 : boolean;
  signal addr_of_1714_final_reg_ack_0 : boolean;
  signal addr_of_1714_final_reg_req_1 : boolean;
  signal type_cast_1832_inst_ack_0 : boolean;
  signal addr_of_1714_final_reg_ack_1 : boolean;
  signal phi_stmt_1829_req_1 : boolean;
  signal type_cast_1834_inst_ack_1 : boolean;
  signal type_cast_1834_inst_req_1 : boolean;
  signal type_cast_1834_inst_ack_0 : boolean;
  signal type_cast_1834_inst_req_0 : boolean;
  signal type_cast_1832_inst_req_0 : boolean;
  signal ptr_deref_1718_load_0_req_0 : boolean;
  signal ptr_deref_1718_load_0_ack_0 : boolean;
  signal phi_stmt_1614_req_0 : boolean;
  signal ptr_deref_1718_load_0_req_1 : boolean;
  signal ptr_deref_1718_load_0_ack_1 : boolean;
  signal phi_stmt_1614_req_1 : boolean;
  signal type_cast_1620_inst_ack_1 : boolean;
  signal type_cast_1620_inst_req_1 : boolean;
  signal type_cast_1620_inst_ack_0 : boolean;
  signal type_cast_1620_inst_req_0 : boolean;
  signal array_obj_ref_1736_index_offset_req_0 : boolean;
  signal array_obj_ref_1736_index_offset_ack_0 : boolean;
  signal array_obj_ref_1736_index_offset_req_1 : boolean;
  signal array_obj_ref_1736_index_offset_ack_1 : boolean;
  signal phi_stmt_1829_ack_0 : boolean;
  signal addr_of_1737_final_reg_req_0 : boolean;
  signal addr_of_1737_final_reg_ack_0 : boolean;
  signal addr_of_1737_final_reg_req_1 : boolean;
  signal addr_of_1737_final_reg_ack_1 : boolean;
  signal ptr_deref_1740_store_0_req_0 : boolean;
  signal ptr_deref_1740_store_0_ack_0 : boolean;
  signal ptr_deref_1740_store_0_req_1 : boolean;
  signal ptr_deref_1740_store_0_ack_1 : boolean;
  signal type_cast_1745_inst_req_0 : boolean;
  signal type_cast_1745_inst_ack_0 : boolean;
  signal type_cast_1745_inst_req_1 : boolean;
  signal type_cast_1745_inst_ack_1 : boolean;
  signal if_stmt_1758_branch_req_0 : boolean;
  signal if_stmt_1758_branch_ack_1 : boolean;
  signal if_stmt_1758_branch_ack_0 : boolean;
  signal type_cast_1786_inst_req_0 : boolean;
  signal type_cast_1786_inst_ack_0 : boolean;
  signal type_cast_1786_inst_req_1 : boolean;
  signal type_cast_1786_inst_ack_1 : boolean;
  signal type_cast_1802_inst_req_0 : boolean;
  signal type_cast_1802_inst_ack_0 : boolean;
  signal type_cast_1802_inst_req_1 : boolean;
  signal type_cast_1802_inst_ack_1 : boolean;
  signal if_stmt_1809_branch_req_0 : boolean;
  signal if_stmt_1809_branch_ack_1 : boolean;
  signal if_stmt_1809_branch_ack_0 : boolean;
  signal WPIPE_Block0_done_1845_inst_req_0 : boolean;
  signal WPIPE_Block0_done_1845_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1845_inst_req_1 : boolean;
  signal WPIPE_Block0_done_1845_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_3763_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3763_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_3763_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3763_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_3763: Block -- control-path 
    signal convTransposeA_CP_3763_elements: BooleanArray(125 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_3763_elements(0) <= convTransposeA_CP_3763_start;
    convTransposeA_CP_3763_symbol <= convTransposeA_CP_3763_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/$entry
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559__entry__
      -- CP-element group 0: 	 branch_block_stmt_1498/$entry
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1498/branch_block_stmt_1498__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_Update/$entry
      -- 
    cr_3956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(0), ack => type_cast_1531_inst_req_1); -- 
    rr_3811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(0), ack => RPIPE_Block0_start_1500_inst_req_0); -- 
    cr_3984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(0), ack => type_cast_1544_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	125 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	84 
    -- CP-element group 1: 	85 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	88 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	91 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	94 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1498/assign_stmt_1841__exit__
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1498/merge_stmt_1815__exit__
      -- CP-element group 1: 	 branch_block_stmt_1498/assign_stmt_1841__entry__
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1628/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/assign_stmt_1841/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/assign_stmt_1841/$exit
      -- 
    cr_4571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(1), ack => type_cast_1634_inst_req_1); -- 
    cr_4502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(1), ack => type_cast_1613_inst_req_1); -- 
    rr_4566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(1), ack => type_cast_1634_inst_req_0); -- 
    cr_4548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(1), ack => type_cast_1627_inst_req_1); -- 
    rr_4497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(1), ack => type_cast_1613_inst_req_0); -- 
    rr_4543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(1), ack => type_cast_1627_inst_req_0); -- 
    cr_4525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(1), ack => type_cast_1620_inst_req_1); -- 
    rr_4520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(1), ack => type_cast_1620_inst_req_0); -- 
    convTransposeA_CP_3763_elements(1) <= convTransposeA_CP_3763_elements(125);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_Update/$entry
      -- 
    ra_3812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1500_inst_ack_0, ack => convTransposeA_CP_3763_elements(2)); -- 
    cr_3816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(2), ack => RPIPE_Block0_start_1500_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_Update/$exit
      -- 
    ca_3817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1500_inst_ack_1, ack => convTransposeA_CP_3763_elements(3)); -- 
    rr_3825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(3), ack => RPIPE_Block0_start_1503_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_Update/$entry
      -- 
    ra_3826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1503_inst_ack_0, ack => convTransposeA_CP_3763_elements(4)); -- 
    cr_3830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(4), ack => RPIPE_Block0_start_1503_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_Update/$exit
      -- 
    ca_3831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1503_inst_ack_1, ack => convTransposeA_CP_3763_elements(5)); -- 
    rr_3839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(5), ack => RPIPE_Block0_start_1506_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_Update/cr
      -- 
    ra_3840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1506_inst_ack_0, ack => convTransposeA_CP_3763_elements(6)); -- 
    cr_3844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(6), ack => RPIPE_Block0_start_1506_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_Sample/rr
      -- 
    ca_3845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1506_inst_ack_1, ack => convTransposeA_CP_3763_elements(7)); -- 
    rr_3853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(7), ack => RPIPE_Block0_start_1509_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_update_start_
      -- 
    ra_3854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1509_inst_ack_0, ack => convTransposeA_CP_3763_elements(8)); -- 
    cr_3858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(8), ack => RPIPE_Block0_start_1509_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_Sample/rr
      -- 
    ca_3859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1509_inst_ack_1, ack => convTransposeA_CP_3763_elements(9)); -- 
    rr_3867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(9), ack => RPIPE_Block0_start_1512_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_Sample/ra
      -- 
    ra_3868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1512_inst_ack_0, ack => convTransposeA_CP_3763_elements(10)); -- 
    cr_3872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(10), ack => RPIPE_Block0_start_1512_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_Update/ca
      -- 
    ca_3873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1512_inst_ack_1, ack => convTransposeA_CP_3763_elements(11)); -- 
    rr_3881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(11), ack => RPIPE_Block0_start_1515_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_Update/cr
      -- 
    ra_3882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1515_inst_ack_0, ack => convTransposeA_CP_3763_elements(12)); -- 
    cr_3886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(12), ack => RPIPE_Block0_start_1515_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_sample_start_
      -- 
    ca_3887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1515_inst_ack_1, ack => convTransposeA_CP_3763_elements(13)); -- 
    rr_3895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(13), ack => RPIPE_Block0_start_1518_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_Update/cr
      -- 
    ra_3896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1518_inst_ack_0, ack => convTransposeA_CP_3763_elements(14)); -- 
    cr_3900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(14), ack => RPIPE_Block0_start_1518_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_Update/ca
      -- 
    ca_3901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1518_inst_ack_1, ack => convTransposeA_CP_3763_elements(15)); -- 
    rr_3909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(15), ack => RPIPE_Block0_start_1521_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_Sample/ra
      -- 
    ra_3910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1521_inst_ack_0, ack => convTransposeA_CP_3763_elements(16)); -- 
    cr_3914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(16), ack => RPIPE_Block0_start_1521_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_Update/ca
      -- 
    ca_3915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1521_inst_ack_1, ack => convTransposeA_CP_3763_elements(17)); -- 
    rr_3923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(17), ack => RPIPE_Block0_start_1524_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_Update/$entry
      -- 
    ra_3924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1524_inst_ack_0, ack => convTransposeA_CP_3763_elements(18)); -- 
    cr_3928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(18), ack => RPIPE_Block0_start_1524_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_Update/$exit
      -- 
    ca_3929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1524_inst_ack_1, ack => convTransposeA_CP_3763_elements(19)); -- 
    rr_3937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(19), ack => RPIPE_Block0_start_1527_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_sample_completed_
      -- 
    ra_3938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1527_inst_ack_0, ack => convTransposeA_CP_3763_elements(20)); -- 
    cr_3942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(20), ack => RPIPE_Block0_start_1527_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_update_completed_
      -- 
    ca_3943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1527_inst_ack_1, ack => convTransposeA_CP_3763_elements(21)); -- 
    rr_3951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(21), ack => type_cast_1531_inst_req_0); -- 
    rr_3965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(21), ack => RPIPE_Block0_start_1540_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_Sample/$exit
      -- 
    ra_3952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1531_inst_ack_0, ack => convTransposeA_CP_3763_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_Update/ca
      -- 
    ca_3957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1531_inst_ack_1, ack => convTransposeA_CP_3763_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_sample_completed_
      -- 
    ra_3966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1540_inst_ack_0, ack => convTransposeA_CP_3763_elements(24)); -- 
    cr_3970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(24), ack => RPIPE_Block0_start_1540_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_Sample/rr
      -- 
    ca_3971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1540_inst_ack_1, ack => convTransposeA_CP_3763_elements(25)); -- 
    rr_3979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(25), ack => type_cast_1544_inst_req_0); -- 
    rr_3993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(25), ack => RPIPE_Block0_start_1552_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_Sample/$exit
      -- 
    ra_3980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1544_inst_ack_0, ack => convTransposeA_CP_3763_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_Update/$exit
      -- 
    ca_3985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1544_inst_ack_1, ack => convTransposeA_CP_3763_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_sample_completed_
      -- 
    ra_3994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1552_inst_ack_0, ack => convTransposeA_CP_3763_elements(28)); -- 
    cr_3998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(28), ack => RPIPE_Block0_start_1552_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_sample_start_
      -- 
    ca_3999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1552_inst_ack_1, ack => convTransposeA_CP_3763_elements(29)); -- 
    rr_4007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(29), ack => RPIPE_Block0_start_1555_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_update_start_
      -- 
    ra_4008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1555_inst_ack_0, ack => convTransposeA_CP_3763_elements(30)); -- 
    cr_4012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(30), ack => RPIPE_Block0_start_1555_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_Sample/rr
      -- 
    ca_4013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1555_inst_ack_1, ack => convTransposeA_CP_3763_elements(31)); -- 
    rr_4021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(31), ack => RPIPE_Block0_start_1558_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_Update/$entry
      -- 
    ra_4022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1558_inst_ack_0, ack => convTransposeA_CP_3763_elements(32)); -- 
    cr_4026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(32), ack => RPIPE_Block0_start_1558_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_update_completed_
      -- 
    ca_4027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1558_inst_ack_1, ack => convTransposeA_CP_3763_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/$exit
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604__entry__
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559__exit__
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1589_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1589_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1589_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1589_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1593_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1593_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1589_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1589_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1585_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1585_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1585_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1585_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1585_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/$entry
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1585_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1593_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1593_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1593_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1593_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1597_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1597_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1597_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1597_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1597_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1597_Update/cr
      -- 
    cr_4057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1589_inst_req_1); -- 
    rr_4052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1589_inst_req_0); -- 
    cr_4043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1585_inst_req_1); -- 
    rr_4038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1585_inst_req_0); -- 
    rr_4066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1593_inst_req_0); -- 
    cr_4071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1593_inst_req_1); -- 
    rr_4080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1597_inst_req_0); -- 
    cr_4085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1597_inst_req_1); -- 
    convTransposeA_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(23) & convTransposeA_CP_3763_elements(27) & convTransposeA_CP_3763_elements(33);
      gj_convTransposeA_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1585_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1585_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1585_sample_completed_
      -- 
    ra_4039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1585_inst_ack_0, ack => convTransposeA_CP_3763_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1585_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1585_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1585_update_completed_
      -- 
    ca_4044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1585_inst_ack_1, ack => convTransposeA_CP_3763_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1589_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1589_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1589_sample_completed_
      -- 
    ra_4053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1589_inst_ack_0, ack => convTransposeA_CP_3763_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1589_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1589_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1589_update_completed_
      -- 
    ca_4058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1589_inst_ack_1, ack => convTransposeA_CP_3763_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1593_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1593_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1593_Sample/ra
      -- 
    ra_4067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1593_inst_ack_0, ack => convTransposeA_CP_3763_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1593_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1593_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1593_Update/ca
      -- 
    ca_4072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1593_inst_ack_1, ack => convTransposeA_CP_3763_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1597_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1597_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1597_Sample/ra
      -- 
    ra_4081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1597_inst_ack_0, ack => convTransposeA_CP_3763_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1597_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1597_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/type_cast_1597_Update/ca
      -- 
    ca_4086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1597_inst_ack_1, ack => convTransposeA_CP_3763_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	82 
    -- CP-element group 43:  members (12) 
      -- CP-element group 43: 	 branch_block_stmt_1498/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604__exit__
      -- CP-element group 43: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1614/$entry
      -- CP-element group 43: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1604/$exit
      -- CP-element group 43: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1621/$entry
      -- CP-element group 43: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1607/$entry
      -- CP-element group 43: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1628/$entry
      -- 
    convTransposeA_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(36) & convTransposeA_CP_3763_elements(38) & convTransposeA_CP_3763_elements(40) & convTransposeA_CP_3763_elements(42);
      gj_convTransposeA_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	102 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1669_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1669_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1669_Sample/ra
      -- 
    ra_4098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1669_inst_ack_0, ack => convTransposeA_CP_3763_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	102 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1669_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1669_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1669_Update/ca
      -- 
    ca_4103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1669_inst_ack_1, ack => convTransposeA_CP_3763_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	102 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1673_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1673_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1673_Sample/ra
      -- 
    ra_4112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1673_inst_ack_0, ack => convTransposeA_CP_3763_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	102 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1673_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1673_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1673_Update/ca
      -- 
    ca_4117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1673_inst_ack_1, ack => convTransposeA_CP_3763_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	102 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1677_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1677_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1677_Sample/ra
      -- 
    ra_4126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1677_inst_ack_0, ack => convTransposeA_CP_3763_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	102 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1677_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1677_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1677_Update/ca
      -- 
    ca_4131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1677_inst_ack_1, ack => convTransposeA_CP_3763_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	102 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1707_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1707_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1707_Sample/ra
      -- 
    ra_4140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1707_inst_ack_0, ack => convTransposeA_CP_3763_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	102 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1707_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1707_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1707_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_final_index_sum_regn_Sample/req
      -- 
    ca_4145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1707_inst_ack_1, ack => convTransposeA_CP_3763_elements(51)); -- 
    req_4170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(51), ack => array_obj_ref_1713_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_final_index_sum_regn_Sample/ack
      -- 
    ack_4171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1713_index_offset_ack_0, ack => convTransposeA_CP_3763_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	102 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1714_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1714_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1714_request/req
      -- 
    ack_4176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1713_index_offset_ack_1, ack => convTransposeA_CP_3763_elements(53)); -- 
    req_4185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(53), ack => addr_of_1714_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1714_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1714_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1714_request/ack
      -- 
    ack_4186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1714_final_reg_ack_0, ack => convTransposeA_CP_3763_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	102 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1714_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1714_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1714_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_Sample/word_access_start/word_0/rr
      -- 
    ack_4191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1714_final_reg_ack_1, ack => convTransposeA_CP_3763_elements(55)); -- 
    rr_4224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(55), ack => ptr_deref_1718_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_Sample/word_access_start/word_0/ra
      -- 
    ra_4225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1718_load_0_ack_0, ack => convTransposeA_CP_3763_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	102 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_Update/ptr_deref_1718_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_Update/ptr_deref_1718_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_Update/ptr_deref_1718_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_Update/ptr_deref_1718_Merge/merge_ack
      -- 
    ca_4236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1718_load_0_ack_1, ack => convTransposeA_CP_3763_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_final_index_sum_regn_Sample/req
      -- 
    req_4266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(58), ack => array_obj_ref_1736_index_offset_req_0); -- 
    convTransposeA_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(45) & convTransposeA_CP_3763_elements(47) & convTransposeA_CP_3763_elements(49);
      gj_convTransposeA_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_final_index_sum_regn_Sample/ack
      -- 
    ack_4267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1736_index_offset_ack_0, ack => convTransposeA_CP_3763_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	102 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1737_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1737_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1737_request/req
      -- 
    ack_4272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1736_index_offset_ack_1, ack => convTransposeA_CP_3763_elements(60)); -- 
    req_4281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(60), ack => addr_of_1737_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1737_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1737_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1737_request/ack
      -- 
    ack_4282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1737_final_reg_ack_0, ack => convTransposeA_CP_3763_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	102 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1737_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1737_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1737_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_word_addrgen/root_register_ack
      -- 
    ack_4287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1737_final_reg_ack_1, ack => convTransposeA_CP_3763_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_Sample/ptr_deref_1740_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_Sample/ptr_deref_1740_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_Sample/ptr_deref_1740_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_Sample/ptr_deref_1740_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_Sample/word_access_start/word_0/rr
      -- 
    rr_4325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(63), ack => ptr_deref_1740_store_0_req_0); -- 
    convTransposeA_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(57) & convTransposeA_CP_3763_elements(62);
      gj_convTransposeA_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_Sample/word_access_start/word_0/ra
      -- 
    ra_4326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1740_store_0_ack_0, ack => convTransposeA_CP_3763_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	102 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_Update/word_access_complete/word_0/ca
      -- 
    ca_4337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1740_store_0_ack_1, ack => convTransposeA_CP_3763_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	102 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1745_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1745_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1745_Sample/ra
      -- 
    ra_4346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1745_inst_ack_0, ack => convTransposeA_CP_3763_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	102 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1745_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1745_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1745_Update/ca
      -- 
    ca_4351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1745_inst_ack_1, ack => convTransposeA_CP_3763_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_1498/if_stmt_1758__entry__
      -- CP-element group 68: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757__exit__
      -- CP-element group 68: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/$exit
      -- CP-element group 68: 	 branch_block_stmt_1498/if_stmt_1758_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1498/if_stmt_1758_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1498/if_stmt_1758_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1498/if_stmt_1758_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1498/R_cmp_1759_place
      -- CP-element group 68: 	 branch_block_stmt_1498/if_stmt_1758_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1498/if_stmt_1758_else_link/$entry
      -- 
    branch_req_4359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(68), ack => if_stmt_1758_branch_req_0); -- 
    convTransposeA_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(52) & convTransposeA_CP_3763_elements(59) & convTransposeA_CP_3763_elements(65) & convTransposeA_CP_3763_elements(67);
      gj_convTransposeA_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	111 
    -- CP-element group 69: 	112 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	115 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	118 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1822/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1498/merge_stmt_1764__exit__
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/assign_stmt_1770__entry__
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1829/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/assign_stmt_1770__exit__
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1822/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123
      -- CP-element group 69: 	 branch_block_stmt_1498/merge_stmt_1764_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1822/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1822/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1822/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1822/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/merge_stmt_1764_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/merge_stmt_1764_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1498/merge_stmt_1764_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1834/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1834/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1834/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1498/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1834/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1834/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1834/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/if_stmt_1758_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1498/if_stmt_1758_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1498/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_1498/assign_stmt_1770/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/assign_stmt_1770/$exit
      -- 
    if_choice_transition_4364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1758_branch_ack_1, ack => convTransposeA_CP_3763_elements(69)); -- 
    cr_4732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(69), ack => type_cast_1822_inst_req_1); -- 
    rr_4727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(69), ack => type_cast_1822_inst_req_0); -- 
    cr_4709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(69), ack => type_cast_1828_inst_req_1); -- 
    rr_4704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(69), ack => type_cast_1828_inst_req_0); -- 
    cr_4686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(69), ack => type_cast_1834_inst_req_1); -- 
    rr_4681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(69), ack => type_cast_1834_inst_req_0); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_1498/merge_stmt_1772_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808__entry__
      -- CP-element group 70: 	 branch_block_stmt_1498/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_1498/merge_stmt_1772_PhiAck/dummy
      -- CP-element group 70: 	 branch_block_stmt_1498/merge_stmt_1772__exit__
      -- CP-element group 70: 	 branch_block_stmt_1498/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1498/merge_stmt_1772_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_1498/merge_stmt_1772_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_1498/if_stmt_1758_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1498/if_stmt_1758_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1498/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/$entry
      -- CP-element group 70: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1786_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1786_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1786_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1786_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1786_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1786_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1802_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1802_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1802_Update/cr
      -- 
    else_choice_transition_4368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1758_branch_ack_0, ack => convTransposeA_CP_3763_elements(70)); -- 
    rr_4384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(70), ack => type_cast_1786_inst_req_0); -- 
    cr_4389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(70), ack => type_cast_1786_inst_req_1); -- 
    cr_4403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(70), ack => type_cast_1802_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1786_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1786_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1786_Sample/ra
      -- 
    ra_4385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1786_inst_ack_0, ack => convTransposeA_CP_3763_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1786_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1786_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1786_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1802_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1802_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1802_Sample/rr
      -- 
    ca_4390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1786_inst_ack_1, ack => convTransposeA_CP_3763_elements(72)); -- 
    rr_4398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(72), ack => type_cast_1802_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1802_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1802_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1802_Sample/ra
      -- 
    ra_4399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1802_inst_ack_0, ack => convTransposeA_CP_3763_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808__exit__
      -- CP-element group 74: 	 branch_block_stmt_1498/if_stmt_1809__entry__
      -- CP-element group 74: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/$exit
      -- CP-element group 74: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1802_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1802_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1498/assign_stmt_1778_to_assign_stmt_1808/type_cast_1802_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_1498/if_stmt_1809_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1498/if_stmt_1809_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1498/if_stmt_1809_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1498/if_stmt_1809_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1498/R_cmp112_1810_place
      -- CP-element group 74: 	 branch_block_stmt_1498/if_stmt_1809_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1498/if_stmt_1809_else_link/$entry
      -- 
    ca_4404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1802_inst_ack_1, ack => convTransposeA_CP_3763_elements(74)); -- 
    branch_req_4412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(74), ack => if_stmt_1809_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_1498/merge_stmt_1843__exit__
      -- CP-element group 75: 	 branch_block_stmt_1498/assign_stmt_1848__entry__
      -- CP-element group 75: 	 branch_block_stmt_1498/merge_stmt_1843_PhiAck/dummy
      -- CP-element group 75: 	 branch_block_stmt_1498/merge_stmt_1843_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1498/merge_stmt_1843_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1498/merge_stmt_1843_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1498/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1498/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1498/if_stmt_1809_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1498/if_stmt_1809_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1498/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_1498/assign_stmt_1848/$entry
      -- CP-element group 75: 	 branch_block_stmt_1498/assign_stmt_1848/WPIPE_Block0_done_1845_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1498/assign_stmt_1848/WPIPE_Block0_done_1845_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1498/assign_stmt_1848/WPIPE_Block0_done_1845_Sample/req
      -- 
    if_choice_transition_4417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1809_branch_ack_1, ack => convTransposeA_CP_3763_elements(75)); -- 
    req_4437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(75), ack => WPIPE_Block0_done_1845_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	103 
    -- CP-element group 76: 	104 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	107 
    -- CP-element group 76: 	109 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1829/$entry
      -- CP-element group 76: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/$entry
      -- CP-element group 76: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/$entry
      -- CP-element group 76: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/$entry
      -- CP-element group 76: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1832/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1832/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1832/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1832/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1832/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1832/$entry
      -- CP-element group 76: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1498/if_stmt_1809_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1498/if_stmt_1809_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123
      -- 
    else_choice_transition_4421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1809_branch_ack_0, ack => convTransposeA_CP_3763_elements(76)); -- 
    cr_4652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(76), ack => type_cast_1826_inst_req_1); -- 
    rr_4647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(76), ack => type_cast_1826_inst_req_0); -- 
    cr_4629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(76), ack => type_cast_1832_inst_req_1); -- 
    rr_4624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(76), ack => type_cast_1832_inst_req_0); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1498/assign_stmt_1848/WPIPE_Block0_done_1845_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1498/assign_stmt_1848/WPIPE_Block0_done_1845_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1498/assign_stmt_1848/WPIPE_Block0_done_1845_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1498/assign_stmt_1848/WPIPE_Block0_done_1845_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1498/assign_stmt_1848/WPIPE_Block0_done_1845_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1498/assign_stmt_1848/WPIPE_Block0_done_1845_Update/req
      -- 
    ack_4438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1845_inst_ack_0, ack => convTransposeA_CP_3763_elements(77)); -- 
    req_4442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(77), ack => WPIPE_Block0_done_1845_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 branch_block_stmt_1498/assign_stmt_1848__exit__
      -- CP-element group 78: 	 branch_block_stmt_1498/return__
      -- CP-element group 78: 	 branch_block_stmt_1498/merge_stmt_1850__exit__
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_1498/$exit
      -- CP-element group 78: 	 branch_block_stmt_1498/merge_stmt_1850_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1498/branch_block_stmt_1498__exit__
      -- CP-element group 78: 	 branch_block_stmt_1498/merge_stmt_1850_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1498/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1498/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1498/merge_stmt_1850_PhiAck/dummy
      -- CP-element group 78: 	 branch_block_stmt_1498/merge_stmt_1850_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1498/assign_stmt_1848/$exit
      -- CP-element group 78: 	 branch_block_stmt_1498/assign_stmt_1848/WPIPE_Block0_done_1845_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1498/assign_stmt_1848/WPIPE_Block0_done_1845_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1498/assign_stmt_1848/WPIPE_Block0_done_1845_Update/ack
      -- 
    ack_4443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1845_inst_ack_1, ack => convTransposeA_CP_3763_elements(78)); -- 
    -- CP-element group 79:  transition  output  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	83 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1611_konst_delay_trans
      -- CP-element group 79: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_req
      -- CP-element group 79: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1607/$exit
      -- 
    phi_stmt_1607_req_4454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1607_req_4454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(79), ack => phi_stmt_1607_req_0); -- 
    -- Element group convTransposeA_CP_3763_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convTransposeA_CP_3763_elements(43), ack => convTransposeA_CP_3763_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  transition  output  delay-element  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1618_konst_delay_trans
      -- CP-element group 80: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1614/$exit
      -- CP-element group 80: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_req
      -- 
    phi_stmt_1614_req_4462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1614_req_4462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(80), ack => phi_stmt_1614_req_0); -- 
    -- Element group convTransposeA_CP_3763_elements(80) is a control-delay.
    cp_element_80_delay: control_delay_element  generic map(name => " 80_delay", delay_value => 1)  port map(req => convTransposeA_CP_3763_elements(43), ack => convTransposeA_CP_3763_elements(80), clk => clk, reset =>reset);
    -- CP-element group 81:  transition  output  delay-element  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	43 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1625_konst_delay_trans
      -- CP-element group 81: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1621/$exit
      -- CP-element group 81: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_req
      -- 
    phi_stmt_1621_req_4470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1621_req_4470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(81), ack => phi_stmt_1621_req_0); -- 
    -- Element group convTransposeA_CP_3763_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => convTransposeA_CP_3763_elements(43), ack => convTransposeA_CP_3763_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  transition  output  delay-element  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1628/phi_stmt_1628_req
      -- CP-element group 82: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1632_konst_delay_trans
      -- CP-element group 82: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/phi_stmt_1628/$exit
      -- 
    phi_stmt_1628_req_4478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1628_req_4478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(82), ack => phi_stmt_1628_req_0); -- 
    -- Element group convTransposeA_CP_3763_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => convTransposeA_CP_3763_elements(43), ack => convTransposeA_CP_3763_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  join  transition  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	79 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	97 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(79) & convTransposeA_CP_3763_elements(80) & convTransposeA_CP_3763_elements(81) & convTransposeA_CP_3763_elements(82);
      gj_convTransposeA_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	1 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/SplitProtocol/Sample/ra
      -- CP-element group 84: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/SplitProtocol/Sample/$exit
      -- 
    ra_4498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1613_inst_ack_0, ack => convTransposeA_CP_3763_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	1 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/SplitProtocol/Update/ca
      -- CP-element group 85: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/SplitProtocol/Update/$exit
      -- 
    ca_4503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1613_inst_ack_1, ack => convTransposeA_CP_3763_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	96 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/$exit
      -- CP-element group 86: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_req
      -- CP-element group 86: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/$exit
      -- CP-element group 86: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/SplitProtocol/$exit
      -- 
    phi_stmt_1607_req_4504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1607_req_4504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(86), ack => phi_stmt_1607_req_1); -- 
    convTransposeA_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(84) & convTransposeA_CP_3763_elements(85);
      gj_convTransposeA_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/SplitProtocol/Sample/ra
      -- CP-element group 87: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/SplitProtocol/Sample/$exit
      -- 
    ra_4521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1620_inst_ack_0, ack => convTransposeA_CP_3763_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	1 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/SplitProtocol/Update/ca
      -- CP-element group 88: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/SplitProtocol/Update/$exit
      -- 
    ca_4526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1620_inst_ack_1, ack => convTransposeA_CP_3763_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	96 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_req
      -- CP-element group 89: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/SplitProtocol/$exit
      -- CP-element group 89: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/$exit
      -- CP-element group 89: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/$exit
      -- 
    phi_stmt_1614_req_4527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1614_req_4527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(89), ack => phi_stmt_1614_req_1); -- 
    convTransposeA_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(87) & convTransposeA_CP_3763_elements(88);
      gj_convTransposeA_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Sample/$exit
      -- 
    ra_4544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1627_inst_ack_0, ack => convTransposeA_CP_3763_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Update/ca
      -- CP-element group 91: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Update/$exit
      -- 
    ca_4549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1627_inst_ack_1, ack => convTransposeA_CP_3763_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	96 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_req
      -- CP-element group 92: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/$exit
      -- CP-element group 92: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/$exit
      -- CP-element group 92: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/$exit
      -- CP-element group 92: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/$exit
      -- 
    phi_stmt_1621_req_4550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1621_req_4550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(92), ack => phi_stmt_1621_req_1); -- 
    convTransposeA_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(90) & convTransposeA_CP_3763_elements(91);
      gj_convTransposeA_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/SplitProtocol/Sample/ra
      -- CP-element group 93: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/SplitProtocol/Sample/$exit
      -- 
    ra_4567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1634_inst_ack_0, ack => convTransposeA_CP_3763_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	1 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/SplitProtocol/Update/ca
      -- CP-element group 94: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/SplitProtocol/Update/$exit
      -- 
    ca_4572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1634_inst_ack_1, ack => convTransposeA_CP_3763_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/$exit
      -- CP-element group 95: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/SplitProtocol/$exit
      -- CP-element group 95: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1628/$exit
      -- CP-element group 95: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1628/phi_stmt_1628_req
      -- CP-element group 95: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/$exit
      -- 
    phi_stmt_1628_req_4573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1628_req_4573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(95), ack => phi_stmt_1628_req_1); -- 
    convTransposeA_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(93) & convTransposeA_CP_3763_elements(94);
      gj_convTransposeA_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	86 
    -- CP-element group 96: 	89 
    -- CP-element group 96: 	92 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_1498/ifx_xend123_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(86) & convTransposeA_CP_3763_elements(89) & convTransposeA_CP_3763_elements(92) & convTransposeA_CP_3763_elements(95);
      gj_convTransposeA_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  merge  fork  transition  place  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	83 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97: 	99 
    -- CP-element group 97: 	100 
    -- CP-element group 97: 	101 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_1498/merge_stmt_1606_PhiAck/$entry
      -- CP-element group 97: 	 branch_block_stmt_1498/merge_stmt_1606_PhiReqMerge
      -- 
    convTransposeA_CP_3763_elements(97) <= OrReduce(convTransposeA_CP_3763_elements(83) & convTransposeA_CP_3763_elements(96));
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	102 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1498/merge_stmt_1606_PhiAck/phi_stmt_1607_ack
      -- 
    phi_stmt_1607_ack_4578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1607_ack_0, ack => convTransposeA_CP_3763_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1498/merge_stmt_1606_PhiAck/phi_stmt_1614_ack
      -- 
    phi_stmt_1614_ack_4579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1614_ack_0, ack => convTransposeA_CP_3763_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	97 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1498/merge_stmt_1606_PhiAck/phi_stmt_1621_ack
      -- 
    phi_stmt_1621_ack_4580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1621_ack_0, ack => convTransposeA_CP_3763_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	97 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1498/merge_stmt_1606_PhiAck/phi_stmt_1628_ack
      -- 
    phi_stmt_1628_ack_4581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1628_ack_0, ack => convTransposeA_CP_3763_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  place  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	98 
    -- CP-element group 102: 	99 
    -- CP-element group 102: 	100 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	44 
    -- CP-element group 102: 	45 
    -- CP-element group 102: 	46 
    -- CP-element group 102: 	47 
    -- CP-element group 102: 	48 
    -- CP-element group 102: 	49 
    -- CP-element group 102: 	50 
    -- CP-element group 102: 	51 
    -- CP-element group 102: 	53 
    -- CP-element group 102: 	55 
    -- CP-element group 102: 	57 
    -- CP-element group 102: 	60 
    -- CP-element group 102: 	62 
    -- CP-element group 102: 	65 
    -- CP-element group 102: 	66 
    -- CP-element group 102: 	67 
    -- CP-element group 102:  members (56) 
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757__entry__
      -- CP-element group 102: 	 branch_block_stmt_1498/merge_stmt_1606__exit__
      -- CP-element group 102: 	 branch_block_stmt_1498/merge_stmt_1606_PhiAck/$exit
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/$entry
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1669_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1669_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1669_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1669_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1669_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1669_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1673_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1673_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1673_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1673_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1673_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1673_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1677_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1677_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1677_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1677_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1677_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1677_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1707_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1707_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1707_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1707_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1707_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1707_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1714_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_final_index_sum_regn_update_start
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_final_index_sum_regn_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1713_final_index_sum_regn_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1714_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1714_complete/req
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_Update/word_access_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_Update/word_access_complete/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1718_Update/word_access_complete/word_0/cr
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1737_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_final_index_sum_regn_update_start
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_final_index_sum_regn_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/array_obj_ref_1736_final_index_sum_regn_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1737_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/addr_of_1737_complete/req
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_Update/word_access_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_Update/word_access_complete/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/ptr_deref_1740_Update/word_access_complete/word_0/cr
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1745_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1745_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1745_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1745_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1745_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1498/assign_stmt_1641_to_assign_stmt_1757/type_cast_1745_Update/cr
      -- 
    rr_4097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => type_cast_1669_inst_req_0); -- 
    cr_4102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => type_cast_1669_inst_req_1); -- 
    rr_4111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => type_cast_1673_inst_req_0); -- 
    cr_4116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => type_cast_1673_inst_req_1); -- 
    rr_4125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => type_cast_1677_inst_req_0); -- 
    cr_4130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => type_cast_1677_inst_req_1); -- 
    rr_4139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => type_cast_1707_inst_req_0); -- 
    cr_4144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => type_cast_1707_inst_req_1); -- 
    req_4175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => array_obj_ref_1713_index_offset_req_1); -- 
    req_4190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => addr_of_1714_final_reg_req_1); -- 
    cr_4235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => ptr_deref_1718_load_0_req_1); -- 
    req_4271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => array_obj_ref_1736_index_offset_req_1); -- 
    req_4286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => addr_of_1737_final_reg_req_1); -- 
    cr_4336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => ptr_deref_1740_store_0_req_1); -- 
    rr_4345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => type_cast_1745_inst_req_0); -- 
    cr_4350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => type_cast_1745_inst_req_1); -- 
    convTransposeA_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(98) & convTransposeA_CP_3763_elements(99) & convTransposeA_CP_3763_elements(100) & convTransposeA_CP_3763_elements(101);
      gj_convTransposeA_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	76 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1832/SplitProtocol/Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1832/SplitProtocol/Sample/$exit
      -- 
    ra_4625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1832_inst_ack_0, ack => convTransposeA_CP_3763_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	76 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1832/SplitProtocol/Update/ca
      -- CP-element group 104: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1832/SplitProtocol/Update/$exit
      -- 
    ca_4630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1832_inst_ack_1, ack => convTransposeA_CP_3763_elements(104)); -- 
    -- CP-element group 105:  join  transition  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	110 
    -- CP-element group 105:  members (5) 
      -- CP-element group 105: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_req
      -- CP-element group 105: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1832/SplitProtocol/$exit
      -- CP-element group 105: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1832/$exit
      -- CP-element group 105: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/$exit
      -- CP-element group 105: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1829/$exit
      -- 
    phi_stmt_1829_req_4631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1829_req_4631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(105), ack => phi_stmt_1829_req_0); -- 
    convTransposeA_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(103) & convTransposeA_CP_3763_elements(104);
      gj_convTransposeA_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Sample/$exit
      -- 
    ra_4648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1826_inst_ack_0, ack => convTransposeA_CP_3763_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	76 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Update/ca
      -- CP-element group 107: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Update/$exit
      -- 
    ca_4653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1826_inst_ack_1, ack => convTransposeA_CP_3763_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_req
      -- CP-element group 108: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/$exit
      -- CP-element group 108: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/$exit
      -- 
    phi_stmt_1823_req_4654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1823_req_4654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(108), ack => phi_stmt_1823_req_0); -- 
    convTransposeA_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(106) & convTransposeA_CP_3763_elements(107);
      gj_convTransposeA_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  output  delay-element  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (4) 
      -- CP-element group 109: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_req
      -- CP-element group 109: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/$exit
      -- CP-element group 109: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1820_konst_delay_trans
      -- CP-element group 109: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/$exit
      -- 
    phi_stmt_1816_req_4662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1816_req_4662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(109), ack => phi_stmt_1816_req_0); -- 
    -- Element group convTransposeA_CP_3763_elements(109) is a control-delay.
    cp_element_109_delay: control_delay_element  generic map(name => " 109_delay", delay_value => 1)  port map(req => convTransposeA_CP_3763_elements(76), ack => convTransposeA_CP_3763_elements(109), clk => clk, reset =>reset);
    -- CP-element group 110:  join  transition  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	105 
    -- CP-element group 110: 	108 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	121 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1498/ifx_xelse_ifx_xend123_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(105) & convTransposeA_CP_3763_elements(108) & convTransposeA_CP_3763_elements(109);
      gj_convTransposeA_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	69 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (2) 
      -- CP-element group 111: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1834/SplitProtocol/Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1834/SplitProtocol/Sample/$exit
      -- 
    ra_4682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1834_inst_ack_0, ack => convTransposeA_CP_3763_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	69 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1834/SplitProtocol/Update/ca
      -- CP-element group 112: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1834/SplitProtocol/Update/$exit
      -- 
    ca_4687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1834_inst_ack_1, ack => convTransposeA_CP_3763_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	120 
    -- CP-element group 113:  members (5) 
      -- CP-element group 113: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1829/$exit
      -- CP-element group 113: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_req
      -- CP-element group 113: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1834/SplitProtocol/$exit
      -- CP-element group 113: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1834/$exit
      -- CP-element group 113: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/$exit
      -- 
    phi_stmt_1829_req_4688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1829_req_4688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(113), ack => phi_stmt_1829_req_1); -- 
    convTransposeA_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(111) & convTransposeA_CP_3763_elements(112);
      gj_convTransposeA_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Sample/$exit
      -- 
    ra_4705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1828_inst_ack_0, ack => convTransposeA_CP_3763_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	69 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Update/ca
      -- CP-element group 115: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Update/$exit
      -- 
    ca_4710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1828_inst_ack_1, ack => convTransposeA_CP_3763_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	120 
    -- CP-element group 116:  members (5) 
      -- CP-element group 116: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_req
      -- CP-element group 116: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/$exit
      -- CP-element group 116: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/$exit
      -- CP-element group 116: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/$exit
      -- CP-element group 116: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/$exit
      -- 
    phi_stmt_1823_req_4711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1823_req_4711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(116), ack => phi_stmt_1823_req_1); -- 
    convTransposeA_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(114) & convTransposeA_CP_3763_elements(115);
      gj_convTransposeA_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1822/SplitProtocol/Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1822/SplitProtocol/Sample/ra
      -- 
    ra_4728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1822_inst_ack_0, ack => convTransposeA_CP_3763_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	69 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1822/SplitProtocol/Update/ca
      -- CP-element group 118: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1822/SplitProtocol/Update/$exit
      -- 
    ca_4733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1822_inst_ack_1, ack => convTransposeA_CP_3763_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1822/$exit
      -- CP-element group 119: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1822/SplitProtocol/$exit
      -- CP-element group 119: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/$exit
      -- CP-element group 119: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/$exit
      -- CP-element group 119: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_req
      -- 
    phi_stmt_1816_req_4734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1816_req_4734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(119), ack => phi_stmt_1816_req_1); -- 
    convTransposeA_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(117) & convTransposeA_CP_3763_elements(118);
      gj_convTransposeA_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	113 
    -- CP-element group 120: 	116 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1498/ifx_xthen_ifx_xend123_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(113) & convTransposeA_CP_3763_elements(116) & convTransposeA_CP_3763_elements(119);
      gj_convTransposeA_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  merge  fork  transition  place  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	110 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: 	123 
    -- CP-element group 121: 	124 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_1498/merge_stmt_1815_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_1498/merge_stmt_1815_PhiReqMerge
      -- 
    convTransposeA_CP_3763_elements(121) <= OrReduce(convTransposeA_CP_3763_elements(110) & convTransposeA_CP_3763_elements(120));
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	125 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1498/merge_stmt_1815_PhiAck/phi_stmt_1816_ack
      -- 
    phi_stmt_1816_ack_4739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1816_ack_0, ack => convTransposeA_CP_3763_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1498/merge_stmt_1815_PhiAck/phi_stmt_1823_ack
      -- 
    phi_stmt_1823_ack_4740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1823_ack_0, ack => convTransposeA_CP_3763_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	121 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1498/merge_stmt_1815_PhiAck/phi_stmt_1829_ack
      -- 
    phi_stmt_1829_ack_4741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1829_ack_0, ack => convTransposeA_CP_3763_elements(124)); -- 
    -- CP-element group 125:  join  transition  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	122 
    -- CP-element group 125: 	123 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	1 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1498/merge_stmt_1815_PhiAck/$exit
      -- 
    convTransposeA_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(122) & convTransposeA_CP_3763_elements(123) & convTransposeA_CP_3763_elements(124);
      gj_convTransposeA_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(125), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom81_1735_resized : std_logic_vector(13 downto 0);
    signal R_idxprom81_1735_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1712_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1712_scaled : std_logic_vector(13 downto 0);
    signal add41_1566 : std_logic_vector(15 downto 0);
    signal add54_1577 : std_logic_vector(15 downto 0);
    signal add73_1688 : std_logic_vector(63 downto 0);
    signal add75_1698 : std_logic_vector(63 downto 0);
    signal add86_1752 : std_logic_vector(31 downto 0);
    signal add93_1770 : std_logic_vector(15 downto 0);
    signal add_1550 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_1646 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1713_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1713_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1713_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1713_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1713_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1713_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1736_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1736_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1736_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1736_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1736_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1736_root_address : std_logic_vector(13 downto 0);
    signal arrayidx77_1715 : std_logic_vector(31 downto 0);
    signal arrayidx82_1738 : std_logic_vector(31 downto 0);
    signal call11_1519 : std_logic_vector(15 downto 0);
    signal call13_1522 : std_logic_vector(15 downto 0);
    signal call14_1525 : std_logic_vector(15 downto 0);
    signal call15_1528 : std_logic_vector(15 downto 0);
    signal call16_1541 : std_logic_vector(15 downto 0);
    signal call18_1553 : std_logic_vector(15 downto 0);
    signal call1_1504 : std_logic_vector(15 downto 0);
    signal call20_1556 : std_logic_vector(15 downto 0);
    signal call22_1559 : std_logic_vector(15 downto 0);
    signal call3_1507 : std_logic_vector(15 downto 0);
    signal call5_1510 : std_logic_vector(15 downto 0);
    signal call7_1513 : std_logic_vector(15 downto 0);
    signal call9_1516 : std_logic_vector(15 downto 0);
    signal call_1501 : std_logic_vector(15 downto 0);
    signal cmp101_1783 : std_logic_vector(0 downto 0);
    signal cmp112_1808 : std_logic_vector(0 downto 0);
    signal cmp_1757 : std_logic_vector(0 downto 0);
    signal conv107_1803 : std_logic_vector(31 downto 0);
    signal conv110_1598 : std_logic_vector(31 downto 0);
    signal conv17_1545 : std_logic_vector(31 downto 0);
    signal conv61_1670 : std_logic_vector(63 downto 0);
    signal conv64_1586 : std_logic_vector(63 downto 0);
    signal conv66_1674 : std_logic_vector(63 downto 0);
    signal conv69_1590 : std_logic_vector(63 downto 0);
    signal conv71_1678 : std_logic_vector(63 downto 0);
    signal conv85_1746 : std_logic_vector(31 downto 0);
    signal conv89_1594 : std_logic_vector(31 downto 0);
    signal conv_1532 : std_logic_vector(31 downto 0);
    signal idxprom81_1731 : std_logic_vector(63 downto 0);
    signal idxprom_1708 : std_logic_vector(63 downto 0);
    signal inc105_1787 : std_logic_vector(15 downto 0);
    signal inc105x_xinput_dim0x_x2_1792 : std_logic_vector(15 downto 0);
    signal inc_1778 : std_logic_vector(15 downto 0);
    signal indvar_1607 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_1841 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_1829 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1628 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_1823 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1621 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1799 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_1816 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1614 : std_logic_vector(15 downto 0);
    signal mul50_1661 : std_logic_vector(15 downto 0);
    signal mul72_1683 : std_logic_vector(63 downto 0);
    signal mul74_1693 : std_logic_vector(63 downto 0);
    signal mul_1651 : std_logic_vector(15 downto 0);
    signal ptr_deref_1718_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1718_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1718_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1718_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1718_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1740_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1740_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1740_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1740_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1740_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1740_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1538 : std_logic_vector(31 downto 0);
    signal shr111126_1604 : std_logic_vector(31 downto 0);
    signal shr80_1725 : std_logic_vector(63 downto 0);
    signal shr_1704 : std_logic_vector(31 downto 0);
    signal sub44_1656 : std_logic_vector(15 downto 0);
    signal sub57_1582 : std_logic_vector(15 downto 0);
    signal sub58_1666 : std_logic_vector(15 downto 0);
    signal sub_1571 : std_logic_vector(15 downto 0);
    signal tmp1_1641 : std_logic_vector(31 downto 0);
    signal tmp78_1719 : std_logic_vector(63 downto 0);
    signal type_cast_1536_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1564_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1575_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1602_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1611_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1613_wire : std_logic_vector(31 downto 0);
    signal type_cast_1618_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1620_wire : std_logic_vector(15 downto 0);
    signal type_cast_1625_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1627_wire : std_logic_vector(15 downto 0);
    signal type_cast_1632_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1634_wire : std_logic_vector(15 downto 0);
    signal type_cast_1639_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1702_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1723_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1729_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1750_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1768_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1776_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1796_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1820_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1822_wire : std_logic_vector(15 downto 0);
    signal type_cast_1826_wire : std_logic_vector(15 downto 0);
    signal type_cast_1828_wire : std_logic_vector(15 downto 0);
    signal type_cast_1832_wire : std_logic_vector(15 downto 0);
    signal type_cast_1834_wire : std_logic_vector(15 downto 0);
    signal type_cast_1839_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1847_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_1713_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1713_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1713_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1713_resized_base_address <= "00000000000000";
    array_obj_ref_1736_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1736_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1736_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1736_resized_base_address <= "00000000000000";
    ptr_deref_1718_word_offset_0 <= "00000000000000";
    ptr_deref_1740_word_offset_0 <= "00000000000000";
    type_cast_1536_wire_constant <= "00000000000000000000000000010000";
    type_cast_1564_wire_constant <= "1111111111111111";
    type_cast_1575_wire_constant <= "1111111111111111";
    type_cast_1602_wire_constant <= "00000000000000000000000000000010";
    type_cast_1611_wire_constant <= "00000000000000000000000000000000";
    type_cast_1618_wire_constant <= "0000000000000000";
    type_cast_1625_wire_constant <= "0000000000000000";
    type_cast_1632_wire_constant <= "0000000000000000";
    type_cast_1639_wire_constant <= "00000000000000000000000000000100";
    type_cast_1702_wire_constant <= "00000000000000000000000000000010";
    type_cast_1723_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1729_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_1750_wire_constant <= "00000000000000000000000000000100";
    type_cast_1768_wire_constant <= "0000000000000100";
    type_cast_1776_wire_constant <= "0000000000000001";
    type_cast_1796_wire_constant <= "0000000000000000";
    type_cast_1820_wire_constant <= "0000000000000000";
    type_cast_1839_wire_constant <= "00000000000000000000000000000001";
    type_cast_1847_wire_constant <= "0000000000000001";
    phi_stmt_1607: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1611_wire_constant & type_cast_1613_wire;
      req <= phi_stmt_1607_req_0 & phi_stmt_1607_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1607",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1607_ack_0,
          idata => idata,
          odata => indvar_1607,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1607
    phi_stmt_1614: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1618_wire_constant & type_cast_1620_wire;
      req <= phi_stmt_1614_req_0 & phi_stmt_1614_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1614",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1614_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1614,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1614
    phi_stmt_1621: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1625_wire_constant & type_cast_1627_wire;
      req <= phi_stmt_1621_req_0 & phi_stmt_1621_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1621",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1621_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1621,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1621
    phi_stmt_1628: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1632_wire_constant & type_cast_1634_wire;
      req <= phi_stmt_1628_req_0 & phi_stmt_1628_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1628",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1628_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1628,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1628
    phi_stmt_1816: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1820_wire_constant & type_cast_1822_wire;
      req <= phi_stmt_1816_req_0 & phi_stmt_1816_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1816",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1816_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_1816,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1816
    phi_stmt_1823: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1826_wire & type_cast_1828_wire;
      req <= phi_stmt_1823_req_0 & phi_stmt_1823_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1823",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1823_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_1823,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1823
    phi_stmt_1829: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1832_wire & type_cast_1834_wire;
      req <= phi_stmt_1829_req_0 & phi_stmt_1829_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1829",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1829_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_1829,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1829
    -- flow-through select operator MUX_1798_inst
    input_dim1x_x2_1799 <= type_cast_1796_wire_constant when (cmp101_1783(0) /=  '0') else inc_1778;
    addr_of_1714_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1714_final_reg_req_0;
      addr_of_1714_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1714_final_reg_req_1;
      addr_of_1714_final_reg_ack_1<= rack(0);
      addr_of_1714_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1714_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1713_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx77_1715,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1737_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1737_final_reg_req_0;
      addr_of_1737_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1737_final_reg_req_1;
      addr_of_1737_final_reg_ack_1<= rack(0);
      addr_of_1737_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1737_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1736_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_1738,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1531_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1531_inst_req_0;
      type_cast_1531_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1531_inst_req_1;
      type_cast_1531_inst_ack_1<= rack(0);
      type_cast_1531_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1531_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1528,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1532,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1544_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1544_inst_req_0;
      type_cast_1544_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1544_inst_req_1;
      type_cast_1544_inst_ack_1<= rack(0);
      type_cast_1544_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1544_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1541,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1545,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1585_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1585_inst_req_0;
      type_cast_1585_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1585_inst_req_1;
      type_cast_1585_inst_ack_1<= rack(0);
      type_cast_1585_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1585_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1559,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv64_1586,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1589_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1589_inst_req_0;
      type_cast_1589_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1589_inst_req_1;
      type_cast_1589_inst_ack_1<= rack(0);
      type_cast_1589_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1589_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1556,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_1590,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1593_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1593_inst_req_0;
      type_cast_1593_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1593_inst_req_1;
      type_cast_1593_inst_ack_1<= rack(0);
      type_cast_1593_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1593_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1507,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv89_1594,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1597_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1597_inst_req_0;
      type_cast_1597_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1597_inst_req_1;
      type_cast_1597_inst_ack_1<= rack(0);
      type_cast_1597_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1597_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1501,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv110_1598,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1613_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1613_inst_req_0;
      type_cast_1613_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1613_inst_req_1;
      type_cast_1613_inst_ack_1<= rack(0);
      type_cast_1613_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1613_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1841,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1613_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1620_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1620_inst_req_0;
      type_cast_1620_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1620_inst_req_1;
      type_cast_1620_inst_ack_1<= rack(0);
      type_cast_1620_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1620_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_1816,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1620_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1627_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1627_inst_req_0;
      type_cast_1627_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1627_inst_req_1;
      type_cast_1627_inst_ack_1<= rack(0);
      type_cast_1627_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1627_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_1823,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1627_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1634_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1634_inst_req_0;
      type_cast_1634_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1634_inst_req_1;
      type_cast_1634_inst_ack_1<= rack(0);
      type_cast_1634_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1634_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_1829,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1634_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1669_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1669_inst_req_0;
      type_cast_1669_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1669_inst_req_1;
      type_cast_1669_inst_ack_1<= rack(0);
      type_cast_1669_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1669_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1614,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_1670,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1673_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1673_inst_req_0;
      type_cast_1673_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1673_inst_req_1;
      type_cast_1673_inst_ack_1<= rack(0);
      type_cast_1673_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1673_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub58_1666,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_1674,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1677_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1677_inst_req_0;
      type_cast_1677_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1677_inst_req_1;
      type_cast_1677_inst_ack_1<= rack(0);
      type_cast_1677_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1677_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub44_1656,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_1678,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1707_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1707_inst_req_0;
      type_cast_1707_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1707_inst_req_1;
      type_cast_1707_inst_ack_1<= rack(0);
      type_cast_1707_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1707_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_1704,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1708,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1745_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1745_inst_req_0;
      type_cast_1745_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1745_inst_req_1;
      type_cast_1745_inst_ack_1<= rack(0);
      type_cast_1745_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1745_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1614,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_1746,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1786_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1786_inst_req_0;
      type_cast_1786_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1786_inst_req_1;
      type_cast_1786_inst_ack_1<= rack(0);
      type_cast_1786_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1786_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp101_1783,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc105_1787,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1802_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1802_inst_req_0;
      type_cast_1802_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1802_inst_req_1;
      type_cast_1802_inst_ack_1<= rack(0);
      type_cast_1802_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1802_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc105x_xinput_dim0x_x2_1792,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_1803,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1822_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1822_inst_req_0;
      type_cast_1822_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1822_inst_req_1;
      type_cast_1822_inst_ack_1<= rack(0);
      type_cast_1822_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1822_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add93_1770,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1822_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1826_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1826_inst_req_0;
      type_cast_1826_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1826_inst_req_1;
      type_cast_1826_inst_ack_1<= rack(0);
      type_cast_1826_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1826_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1799,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1826_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1828_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1828_inst_req_0;
      type_cast_1828_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1828_inst_req_1;
      type_cast_1828_inst_ack_1<= rack(0);
      type_cast_1828_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1828_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1621,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1828_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1832_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1832_inst_req_0;
      type_cast_1832_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1832_inst_req_1;
      type_cast_1832_inst_ack_1<= rack(0);
      type_cast_1832_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1832_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc105x_xinput_dim0x_x2_1792,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1832_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1834_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1834_inst_req_0;
      type_cast_1834_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1834_inst_req_1;
      type_cast_1834_inst_ack_1<= rack(0);
      type_cast_1834_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1834_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1628,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1834_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1713_index_1_rename
    process(R_idxprom_1712_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1712_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1712_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1713_index_1_resize
    process(idxprom_1708) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1708;
      ov := iv(13 downto 0);
      R_idxprom_1712_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1713_root_address_inst
    process(array_obj_ref_1713_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1713_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1713_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1736_index_1_rename
    process(R_idxprom81_1735_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom81_1735_resized;
      ov(13 downto 0) := iv;
      R_idxprom81_1735_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1736_index_1_resize
    process(idxprom81_1731) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom81_1731;
      ov := iv(13 downto 0);
      R_idxprom81_1735_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1736_root_address_inst
    process(array_obj_ref_1736_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1736_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1736_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1718_addr_0
    process(ptr_deref_1718_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1718_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1718_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1718_base_resize
    process(arrayidx77_1715) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx77_1715;
      ov := iv(13 downto 0);
      ptr_deref_1718_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1718_gather_scatter
    process(ptr_deref_1718_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1718_data_0;
      ov(63 downto 0) := iv;
      tmp78_1719 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1718_root_address_inst
    process(ptr_deref_1718_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1718_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1718_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1740_addr_0
    process(ptr_deref_1740_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1740_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1740_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1740_base_resize
    process(arrayidx82_1738) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_1738;
      ov := iv(13 downto 0);
      ptr_deref_1740_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1740_gather_scatter
    process(tmp78_1719) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp78_1719;
      ov(63 downto 0) := iv;
      ptr_deref_1740_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1740_root_address_inst
    process(ptr_deref_1740_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1740_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1740_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1758_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1757;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1758_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1758_branch_req_0,
          ack0 => if_stmt_1758_branch_ack_0,
          ack1 => if_stmt_1758_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1809_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp112_1808;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1809_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1809_branch_req_0,
          ack0 => if_stmt_1809_branch_ack_0,
          ack1 => if_stmt_1809_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1565_inst
    process(call7_1513) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1513, type_cast_1564_wire_constant, tmp_var);
      add41_1566 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1576_inst
    process(call9_1516) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1516, type_cast_1575_wire_constant, tmp_var);
      add54_1577 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1655_inst
    process(sub_1571, mul_1651) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1571, mul_1651, tmp_var);
      sub44_1656 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1665_inst
    process(sub57_1582, mul50_1661) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub57_1582, mul50_1661, tmp_var);
      sub58_1666 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1769_inst
    process(input_dim2x_x1_1614) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1614, type_cast_1768_wire_constant, tmp_var);
      add93_1770 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1777_inst
    process(input_dim1x_x1_1621) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1621, type_cast_1776_wire_constant, tmp_var);
      inc_1778 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1791_inst
    process(inc105_1787, input_dim0x_x2_1628) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc105_1787, input_dim0x_x2_1628, tmp_var);
      inc105x_xinput_dim0x_x2_1792 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1645_inst
    process(add_1550, tmp1_1641) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1550, tmp1_1641, tmp_var);
      add_src_0x_x0_1646 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1751_inst
    process(conv85_1746) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv85_1746, type_cast_1750_wire_constant, tmp_var);
      add86_1752 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1840_inst
    process(indvar_1607) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1607, type_cast_1839_wire_constant, tmp_var);
      indvarx_xnext_1841 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1687_inst
    process(mul72_1683, conv66_1674) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul72_1683, conv66_1674, tmp_var);
      add73_1688 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1697_inst
    process(mul74_1693, conv61_1670) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul74_1693, conv61_1670, tmp_var);
      add75_1698 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1730_inst
    process(shr80_1725) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr80_1725, type_cast_1729_wire_constant, tmp_var);
      idxprom81_1731 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1782_inst
    process(inc_1778, call1_1504) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_1778, call1_1504, tmp_var);
      cmp101_1783 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1807_inst
    process(conv107_1803, shr111126_1604) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv107_1803, shr111126_1604, tmp_var);
      cmp112_1808 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1603_inst
    process(conv110_1598) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv110_1598, type_cast_1602_wire_constant, tmp_var);
      shr111126_1604 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1703_inst
    process(add_src_0x_x0_1646) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_1646, type_cast_1702_wire_constant, tmp_var);
      shr_1704 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1724_inst
    process(add75_1698) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add75_1698, type_cast_1723_wire_constant, tmp_var);
      shr80_1725 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1650_inst
    process(input_dim0x_x2_1628, call13_1522) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_1628, call13_1522, tmp_var);
      mul_1651 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1660_inst
    process(input_dim1x_x1_1621, call13_1522) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1621, call13_1522, tmp_var);
      mul50_1661 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1640_inst
    process(indvar_1607) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1607, type_cast_1639_wire_constant, tmp_var);
      tmp1_1641 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1682_inst
    process(conv71_1678, conv69_1590) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv71_1678, conv69_1590, tmp_var);
      mul72_1683 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1692_inst
    process(add73_1688, conv64_1586) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_1688, conv64_1586, tmp_var);
      mul74_1693 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1549_inst
    process(shl_1538, conv17_1545) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1538, conv17_1545, tmp_var);
      add_1550 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1537_inst
    process(conv_1532) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1532, type_cast_1536_wire_constant, tmp_var);
      shl_1538 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1570_inst
    process(add41_1566, call14_1525) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add41_1566, call14_1525, tmp_var);
      sub_1571 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1581_inst
    process(add54_1577, call14_1525) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add54_1577, call14_1525, tmp_var);
      sub57_1582 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1756_inst
    process(add86_1752, conv89_1594) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add86_1752, conv89_1594, tmp_var);
      cmp_1757 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_1713_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1712_scaled;
      array_obj_ref_1713_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1713_index_offset_req_0;
      array_obj_ref_1713_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1713_index_offset_req_1;
      array_obj_ref_1713_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_1736_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom81_1735_scaled;
      array_obj_ref_1736_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1736_index_offset_req_0;
      array_obj_ref_1736_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1736_index_offset_req_1;
      array_obj_ref_1736_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared load operator group (0) : ptr_deref_1718_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1718_load_0_req_0;
      ptr_deref_1718_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1718_load_0_req_1;
      ptr_deref_1718_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1718_word_address_0;
      ptr_deref_1718_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1740_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1740_store_0_req_0;
      ptr_deref_1740_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1740_store_0_req_1;
      ptr_deref_1740_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1740_word_address_0;
      data_in <= ptr_deref_1740_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1509_inst RPIPE_Block0_start_1515_inst RPIPE_Block0_start_1512_inst RPIPE_Block0_start_1506_inst RPIPE_Block0_start_1503_inst RPIPE_Block0_start_1500_inst RPIPE_Block0_start_1558_inst RPIPE_Block0_start_1555_inst RPIPE_Block0_start_1552_inst RPIPE_Block0_start_1540_inst RPIPE_Block0_start_1527_inst RPIPE_Block0_start_1524_inst RPIPE_Block0_start_1521_inst RPIPE_Block0_start_1518_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block0_start_1509_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block0_start_1515_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block0_start_1512_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block0_start_1506_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block0_start_1503_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block0_start_1500_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block0_start_1558_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block0_start_1555_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block0_start_1552_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block0_start_1540_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block0_start_1527_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block0_start_1524_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block0_start_1521_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block0_start_1518_inst_req_0;
      RPIPE_Block0_start_1509_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block0_start_1515_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block0_start_1512_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block0_start_1506_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block0_start_1503_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block0_start_1500_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block0_start_1558_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block0_start_1555_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block0_start_1552_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block0_start_1540_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block0_start_1527_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block0_start_1524_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block0_start_1521_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block0_start_1518_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block0_start_1509_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block0_start_1515_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block0_start_1512_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block0_start_1506_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block0_start_1503_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block0_start_1500_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block0_start_1558_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block0_start_1555_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block0_start_1552_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block0_start_1540_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block0_start_1527_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block0_start_1524_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block0_start_1521_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block0_start_1518_inst_req_1;
      RPIPE_Block0_start_1509_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block0_start_1515_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block0_start_1512_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block0_start_1506_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block0_start_1503_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block0_start_1500_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block0_start_1558_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block0_start_1555_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block0_start_1552_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block0_start_1540_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block0_start_1527_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block0_start_1524_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block0_start_1521_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block0_start_1518_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call5_1510 <= data_out(223 downto 208);
      call9_1516 <= data_out(207 downto 192);
      call7_1513 <= data_out(191 downto 176);
      call3_1507 <= data_out(175 downto 160);
      call1_1504 <= data_out(159 downto 144);
      call_1501 <= data_out(143 downto 128);
      call22_1559 <= data_out(127 downto 112);
      call20_1556 <= data_out(111 downto 96);
      call18_1553 <= data_out(95 downto 80);
      call16_1541 <= data_out(79 downto 64);
      call15_1528 <= data_out(63 downto 48);
      call14_1525 <= data_out(47 downto 32);
      call13_1522 <= data_out(31 downto 16);
      call11_1519 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1845_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1845_inst_req_0;
      WPIPE_Block0_done_1845_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1845_inst_req_1;
      WPIPE_Block0_done_1845_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1847_wire_constant;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_4758_start: Boolean;
  signal convTransposeB_CP_4758_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block1_start_1862_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1871_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1871_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1868_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1868_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1874_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1874_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1874_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1874_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1862_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1868_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1856_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1856_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1856_inst_req_1 : boolean;
  signal type_cast_1900_inst_ack_1 : boolean;
  signal type_cast_1900_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1908_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1880_inst_req_0 : boolean;
  signal type_cast_1887_inst_ack_0 : boolean;
  signal type_cast_1887_inst_req_0 : boolean;
  signal type_cast_1947_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1883_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1914_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1914_inst_ack_0 : boolean;
  signal type_cast_2189_inst_req_0 : boolean;
  signal type_cast_1900_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1883_inst_req_0 : boolean;
  signal type_cast_2189_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1880_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1862_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1880_inst_req_1 : boolean;
  signal type_cast_1900_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1914_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1914_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1908_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1880_inst_ack_0 : boolean;
  signal type_cast_1947_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1908_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1856_inst_ack_1 : boolean;
  signal type_cast_2193_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1908_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1896_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1865_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1865_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1862_inst_req_0 : boolean;
  signal phi_stmt_2177_req_1 : boolean;
  signal type_cast_2030_inst_req_0 : boolean;
  signal type_cast_2030_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1896_inst_req_1 : boolean;
  signal type_cast_1959_inst_ack_1 : boolean;
  signal type_cast_1959_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1896_inst_ack_0 : boolean;
  signal type_cast_1959_inst_req_0 : boolean;
  signal type_cast_1959_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1896_inst_req_0 : boolean;
  signal phi_stmt_2184_ack_0 : boolean;
  signal RPIPE_Block1_start_1877_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1877_inst_req_1 : boolean;
  signal type_cast_1951_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1871_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1865_inst_ack_0 : boolean;
  signal type_cast_1955_inst_req_0 : boolean;
  signal type_cast_1955_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1871_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1865_inst_req_0 : boolean;
  signal type_cast_1955_inst_req_1 : boolean;
  signal type_cast_1955_inst_ack_1 : boolean;
  signal type_cast_1887_inst_ack_1 : boolean;
  signal type_cast_1887_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1877_inst_ack_0 : boolean;
  signal phi_stmt_2177_ack_0 : boolean;
  signal RPIPE_Block1_start_1877_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1859_inst_ack_1 : boolean;
  signal phi_stmt_2190_ack_0 : boolean;
  signal RPIPE_Block1_start_1859_inst_req_1 : boolean;
  signal type_cast_1951_inst_ack_1 : boolean;
  signal type_cast_1951_inst_req_1 : boolean;
  signal type_cast_2030_inst_req_1 : boolean;
  signal type_cast_2030_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1859_inst_ack_0 : boolean;
  signal type_cast_1947_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1859_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1911_inst_ack_0 : boolean;
  signal type_cast_2189_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1883_inst_ack_1 : boolean;
  signal type_cast_1947_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1883_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1868_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1911_inst_req_0 : boolean;
  signal type_cast_1951_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1911_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1911_inst_ack_1 : boolean;
  signal type_cast_2193_inst_ack_0 : boolean;
  signal type_cast_2034_inst_req_0 : boolean;
  signal type_cast_2034_inst_ack_0 : boolean;
  signal type_cast_2034_inst_req_1 : boolean;
  signal type_cast_2034_inst_ack_1 : boolean;
  signal phi_stmt_2184_req_0 : boolean;
  signal type_cast_2038_inst_req_0 : boolean;
  signal type_cast_2038_inst_ack_0 : boolean;
  signal type_cast_2193_inst_req_0 : boolean;
  signal type_cast_2038_inst_req_1 : boolean;
  signal type_cast_2038_inst_ack_1 : boolean;
  signal type_cast_2187_inst_ack_1 : boolean;
  signal type_cast_2068_inst_req_0 : boolean;
  signal type_cast_2068_inst_ack_0 : boolean;
  signal type_cast_2068_inst_req_1 : boolean;
  signal type_cast_2068_inst_ack_1 : boolean;
  signal type_cast_2187_inst_req_1 : boolean;
  signal type_cast_2187_inst_ack_0 : boolean;
  signal type_cast_2187_inst_req_0 : boolean;
  signal array_obj_ref_2074_index_offset_req_0 : boolean;
  signal array_obj_ref_2074_index_offset_ack_0 : boolean;
  signal array_obj_ref_2074_index_offset_req_1 : boolean;
  signal array_obj_ref_2074_index_offset_ack_1 : boolean;
  signal addr_of_2075_final_reg_req_0 : boolean;
  signal addr_of_2075_final_reg_ack_0 : boolean;
  signal addr_of_2075_final_reg_req_1 : boolean;
  signal addr_of_2075_final_reg_ack_1 : boolean;
  signal ptr_deref_2079_load_0_req_0 : boolean;
  signal ptr_deref_2079_load_0_ack_0 : boolean;
  signal ptr_deref_2079_load_0_req_1 : boolean;
  signal ptr_deref_2079_load_0_ack_1 : boolean;
  signal array_obj_ref_2097_index_offset_req_0 : boolean;
  signal array_obj_ref_2097_index_offset_ack_0 : boolean;
  signal array_obj_ref_2097_index_offset_req_1 : boolean;
  signal array_obj_ref_2097_index_offset_ack_1 : boolean;
  signal phi_stmt_2177_req_0 : boolean;
  signal addr_of_2098_final_reg_req_0 : boolean;
  signal addr_of_2098_final_reg_ack_0 : boolean;
  signal addr_of_2098_final_reg_req_1 : boolean;
  signal addr_of_2098_final_reg_ack_1 : boolean;
  signal type_cast_2180_inst_ack_1 : boolean;
  signal type_cast_2180_inst_req_1 : boolean;
  signal ptr_deref_2101_store_0_req_0 : boolean;
  signal ptr_deref_2101_store_0_ack_0 : boolean;
  signal phi_stmt_2190_req_1 : boolean;
  signal ptr_deref_2101_store_0_req_1 : boolean;
  signal type_cast_2180_inst_ack_0 : boolean;
  signal ptr_deref_2101_store_0_ack_1 : boolean;
  signal type_cast_2180_inst_req_0 : boolean;
  signal type_cast_2106_inst_req_0 : boolean;
  signal type_cast_2106_inst_ack_0 : boolean;
  signal type_cast_2106_inst_req_1 : boolean;
  signal type_cast_2106_inst_ack_1 : boolean;
  signal type_cast_2195_inst_ack_1 : boolean;
  signal if_stmt_2119_branch_req_0 : boolean;
  signal type_cast_2195_inst_req_1 : boolean;
  signal if_stmt_2119_branch_ack_1 : boolean;
  signal if_stmt_2119_branch_ack_0 : boolean;
  signal type_cast_2195_inst_ack_0 : boolean;
  signal type_cast_2195_inst_req_0 : boolean;
  signal type_cast_2147_inst_req_0 : boolean;
  signal type_cast_2147_inst_ack_0 : boolean;
  signal type_cast_2147_inst_req_1 : boolean;
  signal type_cast_2147_inst_ack_1 : boolean;
  signal type_cast_2163_inst_req_0 : boolean;
  signal type_cast_2163_inst_ack_0 : boolean;
  signal type_cast_2163_inst_req_1 : boolean;
  signal type_cast_2163_inst_ack_1 : boolean;
  signal if_stmt_2170_branch_req_0 : boolean;
  signal if_stmt_2170_branch_ack_1 : boolean;
  signal if_stmt_2170_branch_ack_0 : boolean;
  signal WPIPE_Block1_done_2206_inst_req_0 : boolean;
  signal WPIPE_Block1_done_2206_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_2206_inst_req_1 : boolean;
  signal WPIPE_Block1_done_2206_inst_ack_1 : boolean;
  signal type_cast_1993_inst_req_0 : boolean;
  signal type_cast_1993_inst_ack_0 : boolean;
  signal type_cast_1993_inst_req_1 : boolean;
  signal type_cast_1993_inst_ack_1 : boolean;
  signal phi_stmt_1990_req_0 : boolean;
  signal phi_stmt_1983_req_1 : boolean;
  signal phi_stmt_1976_req_0 : boolean;
  signal phi_stmt_1969_req_0 : boolean;
  signal type_cast_1995_inst_req_0 : boolean;
  signal type_cast_1995_inst_ack_0 : boolean;
  signal type_cast_1995_inst_req_1 : boolean;
  signal type_cast_1995_inst_ack_1 : boolean;
  signal phi_stmt_1990_req_1 : boolean;
  signal phi_stmt_2184_req_1 : boolean;
  signal type_cast_1986_inst_req_0 : boolean;
  signal type_cast_1986_inst_ack_0 : boolean;
  signal type_cast_1986_inst_req_1 : boolean;
  signal type_cast_1986_inst_ack_1 : boolean;
  signal phi_stmt_1983_req_0 : boolean;
  signal type_cast_2189_inst_ack_1 : boolean;
  signal type_cast_1982_inst_req_0 : boolean;
  signal type_cast_1982_inst_ack_0 : boolean;
  signal phi_stmt_2190_req_0 : boolean;
  signal type_cast_1982_inst_req_1 : boolean;
  signal type_cast_2193_inst_ack_1 : boolean;
  signal type_cast_1982_inst_ack_1 : boolean;
  signal phi_stmt_1976_req_1 : boolean;
  signal type_cast_1975_inst_req_0 : boolean;
  signal type_cast_1975_inst_ack_0 : boolean;
  signal type_cast_1975_inst_req_1 : boolean;
  signal type_cast_1975_inst_ack_1 : boolean;
  signal phi_stmt_1969_req_1 : boolean;
  signal phi_stmt_1969_ack_0 : boolean;
  signal phi_stmt_1976_ack_0 : boolean;
  signal phi_stmt_1983_ack_0 : boolean;
  signal phi_stmt_1990_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_4758_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4758_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_4758_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4758_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_4758: Block -- control-path 
    signal convTransposeB_CP_4758_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_4758_elements(0) <= convTransposeB_CP_4758_start;
    convTransposeB_CP_4758_symbol <= convTransposeB_CP_4758_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_1854/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1854/branch_block_stmt_1854__entry__
      -- CP-element group 0: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915__entry__
      -- CP-element group 0: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1856_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1856_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1900_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1856_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1900_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/$entry
      -- CP-element group 0: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1887_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1900_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1887_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1887_Update/$entry
      -- 
    rr_4806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(0), ack => RPIPE_Block1_start_1856_inst_req_0); -- 
    cr_4979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(0), ack => type_cast_1900_inst_req_1); -- 
    cr_4951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(0), ack => type_cast_1887_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	92 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1854/merge_stmt_2176__exit__
      -- CP-element group 1: 	 branch_block_stmt_1854/assign_stmt_2202__entry__
      -- CP-element group 1: 	 branch_block_stmt_1854/assign_stmt_2202__exit__
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1854/assign_stmt_2202/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/assign_stmt_2202/$exit
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1990/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1995/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1995/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1995/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1995/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1995/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1995/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/SplitProtocol/Update/cr
      -- 
    rr_5507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(1), ack => type_cast_1995_inst_req_0); -- 
    cr_5512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(1), ack => type_cast_1995_inst_req_1); -- 
    rr_5530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(1), ack => type_cast_1986_inst_req_0); -- 
    cr_5535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(1), ack => type_cast_1986_inst_req_1); -- 
    rr_5553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(1), ack => type_cast_1982_inst_req_0); -- 
    cr_5558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(1), ack => type_cast_1982_inst_req_1); -- 
    rr_5576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(1), ack => type_cast_1975_inst_req_0); -- 
    cr_5581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(1), ack => type_cast_1975_inst_req_1); -- 
    convTransposeB_CP_4758_elements(1) <= convTransposeB_CP_4758_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1856_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1856_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1856_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1856_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1856_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1856_sample_completed_
      -- 
    ra_4807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1856_inst_ack_0, ack => convTransposeB_CP_4758_elements(2)); -- 
    cr_4811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(2), ack => RPIPE_Block1_start_1856_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1859_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1856_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1856_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1856_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1859_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1859_Sample/$entry
      -- 
    ca_4812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1856_inst_ack_1, ack => convTransposeB_CP_4758_elements(3)); -- 
    rr_4820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(3), ack => RPIPE_Block1_start_1859_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1859_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1859_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1859_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1859_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1859_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1859_Sample/$exit
      -- 
    ra_4821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1859_inst_ack_0, ack => convTransposeB_CP_4758_elements(4)); -- 
    cr_4825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(4), ack => RPIPE_Block1_start_1859_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1862_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1859_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1862_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1862_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1859_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1859_Update/$exit
      -- 
    ca_4826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1859_inst_ack_1, ack => convTransposeB_CP_4758_elements(5)); -- 
    rr_4834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(5), ack => RPIPE_Block1_start_1862_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1862_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1862_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1862_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1862_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1862_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1862_sample_completed_
      -- 
    ra_4835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1862_inst_ack_0, ack => convTransposeB_CP_4758_elements(6)); -- 
    cr_4839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(6), ack => RPIPE_Block1_start_1862_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1862_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1862_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1865_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1862_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1865_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1865_Sample/$entry
      -- 
    ca_4840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1862_inst_ack_1, ack => convTransposeB_CP_4758_elements(7)); -- 
    rr_4848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(7), ack => RPIPE_Block1_start_1865_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1865_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1865_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1865_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1865_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1865_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1865_update_start_
      -- 
    ra_4849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1865_inst_ack_0, ack => convTransposeB_CP_4758_elements(8)); -- 
    cr_4853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(8), ack => RPIPE_Block1_start_1865_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1868_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1868_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1868_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1865_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1865_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1865_update_completed_
      -- 
    ca_4854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1865_inst_ack_1, ack => convTransposeB_CP_4758_elements(9)); -- 
    rr_4862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(9), ack => RPIPE_Block1_start_1868_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1868_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1868_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1868_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1868_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1868_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1868_Sample/ra
      -- 
    ra_4863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1868_inst_ack_0, ack => convTransposeB_CP_4758_elements(10)); -- 
    cr_4867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(10), ack => RPIPE_Block1_start_1868_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1868_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1871_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1868_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1868_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1871_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1871_Sample/$entry
      -- 
    ca_4868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1868_inst_ack_1, ack => convTransposeB_CP_4758_elements(11)); -- 
    rr_4876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(11), ack => RPIPE_Block1_start_1871_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1871_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1871_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1871_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1871_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1871_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1871_Sample/$exit
      -- 
    ra_4877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1871_inst_ack_0, ack => convTransposeB_CP_4758_elements(12)); -- 
    cr_4881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(12), ack => RPIPE_Block1_start_1871_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1871_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1874_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1874_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1871_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1874_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1871_update_completed_
      -- 
    ca_4882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1871_inst_ack_1, ack => convTransposeB_CP_4758_elements(13)); -- 
    rr_4890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(13), ack => RPIPE_Block1_start_1874_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1874_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1874_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1874_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1874_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1874_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1874_update_start_
      -- 
    ra_4891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1874_inst_ack_0, ack => convTransposeB_CP_4758_elements(14)); -- 
    cr_4895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(14), ack => RPIPE_Block1_start_1874_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1874_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1874_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1877_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1874_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1877_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1877_Sample/$entry
      -- 
    ca_4896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1874_inst_ack_1, ack => convTransposeB_CP_4758_elements(15)); -- 
    rr_4904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(15), ack => RPIPE_Block1_start_1877_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1877_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1877_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1877_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1877_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1877_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1877_Sample/ra
      -- 
    ra_4905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1877_inst_ack_0, ack => convTransposeB_CP_4758_elements(16)); -- 
    cr_4909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(16), ack => RPIPE_Block1_start_1877_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1880_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1880_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1880_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1877_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1877_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1877_update_completed_
      -- 
    ca_4910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1877_inst_ack_1, ack => convTransposeB_CP_4758_elements(17)); -- 
    rr_4918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(17), ack => RPIPE_Block1_start_1880_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1880_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1880_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1880_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1880_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1880_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1880_sample_completed_
      -- 
    ra_4919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1880_inst_ack_0, ack => convTransposeB_CP_4758_elements(18)); -- 
    cr_4923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(18), ack => RPIPE_Block1_start_1880_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1883_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1883_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1880_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1883_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1880_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1880_update_completed_
      -- 
    ca_4924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1880_inst_ack_1, ack => convTransposeB_CP_4758_elements(19)); -- 
    rr_4932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(19), ack => RPIPE_Block1_start_1883_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1883_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1883_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1883_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1883_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1883_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1883_Update/cr
      -- 
    ra_4933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1883_inst_ack_0, ack => convTransposeB_CP_4758_elements(20)); -- 
    cr_4937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(20), ack => RPIPE_Block1_start_1883_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1887_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1883_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1887_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1883_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1896_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1896_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1896_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1887_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1883_Update/ca
      -- 
    ca_4938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1883_inst_ack_1, ack => convTransposeB_CP_4758_elements(21)); -- 
    rr_4946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(21), ack => type_cast_1887_inst_req_0); -- 
    rr_4960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(21), ack => RPIPE_Block1_start_1896_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1887_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1887_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1887_sample_completed_
      -- 
    ra_4947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1887_inst_ack_0, ack => convTransposeB_CP_4758_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1887_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1887_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1887_Update/$exit
      -- 
    ca_4952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1887_inst_ack_1, ack => convTransposeB_CP_4758_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1896_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1896_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1896_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1896_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1896_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1896_sample_completed_
      -- 
    ra_4961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1896_inst_ack_0, ack => convTransposeB_CP_4758_elements(24)); -- 
    cr_4965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(24), ack => RPIPE_Block1_start_1896_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1908_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1900_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1900_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1900_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1908_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1896_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1908_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1896_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1896_update_completed_
      -- 
    ca_4966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1896_inst_ack_1, ack => convTransposeB_CP_4758_elements(25)); -- 
    rr_4974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(25), ack => type_cast_1900_inst_req_0); -- 
    rr_4988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(25), ack => RPIPE_Block1_start_1908_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1900_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1900_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1900_Sample/ra
      -- 
    ra_4975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1900_inst_ack_0, ack => convTransposeB_CP_4758_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1900_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1900_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/type_cast_1900_Update/$exit
      -- 
    ca_4980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1900_inst_ack_1, ack => convTransposeB_CP_4758_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1908_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1908_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1908_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1908_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1908_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1908_Update/$entry
      -- 
    ra_4989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1908_inst_ack_0, ack => convTransposeB_CP_4758_elements(28)); -- 
    cr_4993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(28), ack => RPIPE_Block1_start_1908_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1911_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1908_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1911_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1908_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1908_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1911_Sample/rr
      -- 
    ca_4994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1908_inst_ack_1, ack => convTransposeB_CP_4758_elements(29)); -- 
    rr_5002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(29), ack => RPIPE_Block1_start_1911_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1911_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1911_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1911_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1911_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1911_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1911_Update/cr
      -- 
    ra_5003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1911_inst_ack_0, ack => convTransposeB_CP_4758_elements(30)); -- 
    cr_5007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(30), ack => RPIPE_Block1_start_1911_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1914_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1914_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1911_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1911_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1914_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1911_Update/ca
      -- 
    ca_5008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1911_inst_ack_1, ack => convTransposeB_CP_4758_elements(31)); -- 
    rr_5016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(31), ack => RPIPE_Block1_start_1914_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1914_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1914_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1914_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1914_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1914_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1914_sample_completed_
      -- 
    ra_5017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1914_inst_ack_0, ack => convTransposeB_CP_4758_elements(32)); -- 
    cr_5021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(32), ack => RPIPE_Block1_start_1914_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1914_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1914_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/RPIPE_Block1_start_1914_Update/ca
      -- 
    ca_5022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1914_inst_ack_1, ack => convTransposeB_CP_4758_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966__entry__
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915__exit__
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/$entry
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1947_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1857_to_assign_stmt_1915/$exit
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1947_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1947_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1947_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1959_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1959_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1959_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1959_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1959_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1959_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1951_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1951_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1955_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1955_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1955_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1955_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1955_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1955_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1951_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1951_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1947_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1947_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1951_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1951_update_start_
      -- 
    rr_5033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(34), ack => type_cast_1947_inst_req_0); -- 
    cr_5080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(34), ack => type_cast_1959_inst_req_1); -- 
    rr_5075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(34), ack => type_cast_1959_inst_req_0); -- 
    rr_5047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(34), ack => type_cast_1951_inst_req_0); -- 
    rr_5061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(34), ack => type_cast_1955_inst_req_0); -- 
    cr_5066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(34), ack => type_cast_1955_inst_req_1); -- 
    cr_5052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(34), ack => type_cast_1951_inst_req_1); -- 
    cr_5038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(34), ack => type_cast_1947_inst_req_1); -- 
    convTransposeB_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(23) & convTransposeB_CP_4758_elements(27) & convTransposeB_CP_4758_elements(33);
      gj_convTransposeB_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1947_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1947_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1947_Sample/$exit
      -- 
    ra_5034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1947_inst_ack_0, ack => convTransposeB_CP_4758_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1947_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1947_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1947_Update/$exit
      -- 
    ca_5039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1947_inst_ack_1, ack => convTransposeB_CP_4758_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1951_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1951_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1951_Sample/ra
      -- 
    ra_5048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1951_inst_ack_0, ack => convTransposeB_CP_4758_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1951_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1951_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1951_update_completed_
      -- 
    ca_5053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1951_inst_ack_1, ack => convTransposeB_CP_4758_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1955_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1955_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1955_sample_completed_
      -- 
    ra_5062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1955_inst_ack_0, ack => convTransposeB_CP_4758_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1955_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1955_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1955_update_completed_
      -- 
    ca_5067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1955_inst_ack_1, ack => convTransposeB_CP_4758_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1959_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1959_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1959_sample_completed_
      -- 
    ra_5076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1959_inst_ack_0, ack => convTransposeB_CP_4758_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1959_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1959_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/type_cast_1959_update_completed_
      -- 
    ca_5081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1959_inst_ack_1, ack => convTransposeB_CP_4758_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	82 
    -- CP-element group 43: 	83 
    -- CP-element group 43: 	84 
    -- CP-element group 43:  members (18) 
      -- CP-element group 43: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966__exit__
      -- CP-element group 43: 	 branch_block_stmt_1854/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1854/assign_stmt_1922_to_assign_stmt_1966/$exit
      -- CP-element group 43: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1990/$entry
      -- CP-element group 43: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1993/$entry
      -- CP-element group 43: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1993/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1993/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1993/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1993/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1993/SplitProtocol/Update/cr
      -- CP-element group 43: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1983/$entry
      -- CP-element group 43: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1976/$entry
      -- CP-element group 43: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1969/$entry
      -- CP-element group 43: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/$entry
      -- 
    rr_5457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(43), ack => type_cast_1993_inst_req_0); -- 
    cr_5462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(43), ack => type_cast_1993_inst_req_1); -- 
    convTransposeB_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(36) & convTransposeB_CP_4758_elements(38) & convTransposeB_CP_4758_elements(40) & convTransposeB_CP_4758_elements(42);
      gj_convTransposeB_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	104 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2030_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2030_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2030_Sample/$exit
      -- 
    ra_5093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2030_inst_ack_0, ack => convTransposeB_CP_4758_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	104 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2030_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2030_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2030_Update/ca
      -- 
    ca_5098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2030_inst_ack_1, ack => convTransposeB_CP_4758_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	104 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2034_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2034_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2034_Sample/ra
      -- 
    ra_5107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2034_inst_ack_0, ack => convTransposeB_CP_4758_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	104 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2034_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2034_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2034_Update/ca
      -- 
    ca_5112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2034_inst_ack_1, ack => convTransposeB_CP_4758_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	104 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2038_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2038_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2038_Sample/ra
      -- 
    ra_5121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2038_inst_ack_0, ack => convTransposeB_CP_4758_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	104 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2038_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2038_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2038_Update/ca
      -- 
    ca_5126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2038_inst_ack_1, ack => convTransposeB_CP_4758_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	104 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2068_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2068_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2068_Sample/ra
      -- 
    ra_5135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2068_inst_ack_0, ack => convTransposeB_CP_4758_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	104 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2068_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2068_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2068_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_final_index_sum_regn_Sample/req
      -- 
    ca_5140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2068_inst_ack_1, ack => convTransposeB_CP_4758_elements(51)); -- 
    req_5165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(51), ack => array_obj_ref_2074_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_final_index_sum_regn_Sample/ack
      -- 
    ack_5166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2074_index_offset_ack_0, ack => convTransposeB_CP_4758_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	104 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2075_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2075_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2075_request/req
      -- 
    ack_5171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2074_index_offset_ack_1, ack => convTransposeB_CP_4758_elements(53)); -- 
    req_5180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(53), ack => addr_of_2075_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2075_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2075_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2075_request/ack
      -- 
    ack_5181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2075_final_reg_ack_0, ack => convTransposeB_CP_4758_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	104 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2075_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2075_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2075_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_Sample/word_access_start/word_0/rr
      -- 
    ack_5186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2075_final_reg_ack_1, ack => convTransposeB_CP_4758_elements(55)); -- 
    rr_5219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(55), ack => ptr_deref_2079_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_Sample/word_access_start/word_0/ra
      -- 
    ra_5220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2079_load_0_ack_0, ack => convTransposeB_CP_4758_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	104 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_Update/ptr_deref_2079_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_Update/ptr_deref_2079_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_Update/ptr_deref_2079_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_Update/ptr_deref_2079_Merge/merge_ack
      -- 
    ca_5231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2079_load_0_ack_1, ack => convTransposeB_CP_4758_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_final_index_sum_regn_Sample/req
      -- 
    req_5261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(58), ack => array_obj_ref_2097_index_offset_req_0); -- 
    convTransposeB_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(45) & convTransposeB_CP_4758_elements(47) & convTransposeB_CP_4758_elements(49);
      gj_convTransposeB_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_final_index_sum_regn_Sample/ack
      -- 
    ack_5262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2097_index_offset_ack_0, ack => convTransposeB_CP_4758_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	104 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2098_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2098_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2098_request/req
      -- 
    ack_5267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2097_index_offset_ack_1, ack => convTransposeB_CP_4758_elements(60)); -- 
    req_5276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(60), ack => addr_of_2098_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2098_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2098_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2098_request/ack
      -- 
    ack_5277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2098_final_reg_ack_0, ack => convTransposeB_CP_4758_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	104 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2098_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2098_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2098_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_word_addrgen/root_register_ack
      -- 
    ack_5282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2098_final_reg_ack_1, ack => convTransposeB_CP_4758_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_Sample/ptr_deref_2101_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_Sample/ptr_deref_2101_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_Sample/ptr_deref_2101_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_Sample/ptr_deref_2101_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_Sample/word_access_start/word_0/rr
      -- 
    rr_5320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(63), ack => ptr_deref_2101_store_0_req_0); -- 
    convTransposeB_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(57) & convTransposeB_CP_4758_elements(62);
      gj_convTransposeB_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_Sample/word_access_start/word_0/ra
      -- 
    ra_5321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2101_store_0_ack_0, ack => convTransposeB_CP_4758_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	104 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_Update/word_access_complete/word_0/ca
      -- 
    ca_5332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2101_store_0_ack_1, ack => convTransposeB_CP_4758_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	104 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2106_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2106_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2106_Sample/ra
      -- 
    ra_5341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2106_inst_ack_0, ack => convTransposeB_CP_4758_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	104 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2106_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2106_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2106_Update/ca
      -- 
    ca_5346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2106_inst_ack_1, ack => convTransposeB_CP_4758_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_1854/if_stmt_2119__entry__
      -- CP-element group 68: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118__exit__
      -- CP-element group 68: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/$exit
      -- CP-element group 68: 	 branch_block_stmt_1854/if_stmt_2119_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1854/if_stmt_2119_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1854/if_stmt_2119_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1854/if_stmt_2119_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1854/R_cmp_2120_place
      -- CP-element group 68: 	 branch_block_stmt_1854/if_stmt_2119_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1854/if_stmt_2119_else_link/$entry
      -- 
    branch_req_5354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(68), ack => if_stmt_2119_branch_req_0); -- 
    convTransposeB_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(52) & convTransposeB_CP_4758_elements(59) & convTransposeB_CP_4758_elements(65) & convTransposeB_CP_4758_elements(67);
      gj_convTransposeB_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	113 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	116 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	119 
    -- CP-element group 69: 	120 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_1854/merge_stmt_2125__exit__
      -- CP-element group 69: 	 branch_block_stmt_1854/assign_stmt_2131__entry__
      -- CP-element group 69: 	 branch_block_stmt_1854/assign_stmt_2131__exit__
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1854/if_stmt_2119_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1854/if_stmt_2119_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1854/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_1854/assign_stmt_2131/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/assign_stmt_2131/$exit
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2190/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1854/merge_stmt_2125_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1854/merge_stmt_2125_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1854/merge_stmt_2125_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1854/merge_stmt_2125_PhiAck/dummy
      -- 
    if_choice_transition_5359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2119_branch_ack_1, ack => convTransposeB_CP_4758_elements(69)); -- 
    cr_5696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(69), ack => type_cast_2193_inst_req_1); -- 
    rr_5691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(69), ack => type_cast_2193_inst_req_0); -- 
    cr_5742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(69), ack => type_cast_2187_inst_req_1); -- 
    rr_5737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(69), ack => type_cast_2187_inst_req_0); -- 
    cr_5719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(69), ack => type_cast_2180_inst_req_1); -- 
    rr_5714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(69), ack => type_cast_2180_inst_req_0); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_1854/merge_stmt_2133__exit__
      -- CP-element group 70: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169__entry__
      -- CP-element group 70: 	 branch_block_stmt_1854/if_stmt_2119_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1854/if_stmt_2119_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1854/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/$entry
      -- CP-element group 70: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2147_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2147_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2147_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2147_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2147_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2147_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2163_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2163_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2163_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1854/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1854/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_1854/merge_stmt_2133_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_1854/merge_stmt_2133_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_1854/merge_stmt_2133_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_1854/merge_stmt_2133_PhiAck/dummy
      -- 
    else_choice_transition_5363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2119_branch_ack_0, ack => convTransposeB_CP_4758_elements(70)); -- 
    rr_5379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(70), ack => type_cast_2147_inst_req_0); -- 
    cr_5384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(70), ack => type_cast_2147_inst_req_1); -- 
    cr_5398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(70), ack => type_cast_2163_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2147_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2147_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2147_Sample/ra
      -- 
    ra_5380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2147_inst_ack_0, ack => convTransposeB_CP_4758_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2147_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2147_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2147_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2163_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2163_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2163_Sample/rr
      -- 
    ca_5385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2147_inst_ack_1, ack => convTransposeB_CP_4758_elements(72)); -- 
    rr_5393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(72), ack => type_cast_2163_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2163_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2163_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2163_Sample/ra
      -- 
    ra_5394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2163_inst_ack_0, ack => convTransposeB_CP_4758_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_1854/if_stmt_2170__entry__
      -- CP-element group 74: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169__exit__
      -- CP-element group 74: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/$exit
      -- CP-element group 74: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2163_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2163_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1854/assign_stmt_2139_to_assign_stmt_2169/type_cast_2163_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_1854/if_stmt_2170_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1854/if_stmt_2170_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1854/if_stmt_2170_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1854/if_stmt_2170_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1854/R_cmp117_2171_place
      -- CP-element group 74: 	 branch_block_stmt_1854/if_stmt_2170_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1854/if_stmt_2170_else_link/$entry
      -- 
    ca_5399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2163_inst_ack_1, ack => convTransposeB_CP_4758_elements(74)); -- 
    branch_req_5407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(74), ack => if_stmt_2170_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_1854/assign_stmt_2209__entry__
      -- CP-element group 75: 	 branch_block_stmt_1854/merge_stmt_2204__exit__
      -- CP-element group 75: 	 branch_block_stmt_1854/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1854/merge_stmt_2204_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1854/merge_stmt_2204_PhiAck/dummy
      -- CP-element group 75: 	 branch_block_stmt_1854/merge_stmt_2204_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1854/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1854/merge_stmt_2204_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1854/if_stmt_2170_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1854/if_stmt_2170_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1854/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_1854/assign_stmt_2209/$entry
      -- CP-element group 75: 	 branch_block_stmt_1854/assign_stmt_2209/WPIPE_Block1_done_2206_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1854/assign_stmt_2209/WPIPE_Block1_done_2206_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1854/assign_stmt_2209/WPIPE_Block1_done_2206_Sample/req
      -- 
    if_choice_transition_5412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2170_branch_ack_1, ack => convTransposeB_CP_4758_elements(75)); -- 
    req_5432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(75), ack => WPIPE_Block1_done_2206_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	105 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	108 
    -- CP-element group 76: 	109 
    -- CP-element group 76: 	110 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/$entry
      -- CP-element group 76: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/$entry
      -- CP-element group 76: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2195/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2195/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2195/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2190/$entry
      -- CP-element group 76: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2195/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1854/if_stmt_2170_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2195/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1854/if_stmt_2170_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128
      -- CP-element group 76: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2195/$entry
      -- CP-element group 76: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/$entry
      -- CP-element group 76: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/$entry
      -- 
    else_choice_transition_5416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2170_branch_ack_0, ack => convTransposeB_CP_4758_elements(76)); -- 
    rr_5665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(76), ack => type_cast_2189_inst_req_0); -- 
    cr_5670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(76), ack => type_cast_2189_inst_req_1); -- 
    cr_5639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(76), ack => type_cast_2195_inst_req_1); -- 
    rr_5634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(76), ack => type_cast_2195_inst_req_0); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1854/assign_stmt_2209/WPIPE_Block1_done_2206_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1854/assign_stmt_2209/WPIPE_Block1_done_2206_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1854/assign_stmt_2209/WPIPE_Block1_done_2206_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1854/assign_stmt_2209/WPIPE_Block1_done_2206_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1854/assign_stmt_2209/WPIPE_Block1_done_2206_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1854/assign_stmt_2209/WPIPE_Block1_done_2206_Update/req
      -- 
    ack_5433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2206_inst_ack_0, ack => convTransposeB_CP_4758_elements(77)); -- 
    req_5437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(77), ack => WPIPE_Block1_done_2206_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_1854/branch_block_stmt_1854__exit__
      -- CP-element group 78: 	 branch_block_stmt_1854/$exit
      -- CP-element group 78: 	 branch_block_stmt_1854/assign_stmt_2209__exit__
      -- CP-element group 78: 	 branch_block_stmt_1854/merge_stmt_2211__exit__
      -- CP-element group 78: 	 branch_block_stmt_1854/return__
      -- CP-element group 78: 	 branch_block_stmt_1854/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1854/merge_stmt_2211_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1854/merge_stmt_2211_PhiAck/dummy
      -- CP-element group 78: 	 branch_block_stmt_1854/merge_stmt_2211_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1854/assign_stmt_2209/$exit
      -- CP-element group 78: 	 branch_block_stmt_1854/assign_stmt_2209/WPIPE_Block1_done_2206_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1854/merge_stmt_2211_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1854/assign_stmt_2209/WPIPE_Block1_done_2206_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1854/assign_stmt_2209/WPIPE_Block1_done_2206_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_1854/return___PhiReq/$exit
      -- 
    ack_5438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2206_inst_ack_1, ack => convTransposeB_CP_4758_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1993/SplitProtocol/Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1993/SplitProtocol/Sample/ra
      -- 
    ra_5458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1993_inst_ack_0, ack => convTransposeB_CP_4758_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1993/SplitProtocol/Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1993/SplitProtocol/Update/ca
      -- 
    ca_5463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1993_inst_ack_1, ack => convTransposeB_CP_4758_elements(80)); -- 
    -- CP-element group 81:  join  transition  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1990/$exit
      -- CP-element group 81: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1993/$exit
      -- CP-element group 81: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1993/SplitProtocol/$exit
      -- CP-element group 81: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_req
      -- 
    phi_stmt_1990_req_5464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1990_req_5464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(81), ack => phi_stmt_1990_req_0); -- 
    convTransposeB_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(79) & convTransposeB_CP_4758_elements(80);
      gj_convTransposeB_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  output  delay-element  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	85 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1983/$exit
      -- CP-element group 82: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1989_konst_delay_trans
      -- CP-element group 82: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_req
      -- 
    phi_stmt_1983_req_5472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1983_req_5472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(82), ack => phi_stmt_1983_req_1); -- 
    -- Element group convTransposeB_CP_4758_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => convTransposeB_CP_4758_elements(43), ack => convTransposeB_CP_4758_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  transition  output  delay-element  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	43 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1976/$exit
      -- CP-element group 83: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/$exit
      -- CP-element group 83: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1980_konst_delay_trans
      -- CP-element group 83: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_req
      -- 
    phi_stmt_1976_req_5480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1976_req_5480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(83), ack => phi_stmt_1976_req_0); -- 
    -- Element group convTransposeB_CP_4758_elements(83) is a control-delay.
    cp_element_83_delay: control_delay_element  generic map(name => " 83_delay", delay_value => 1)  port map(req => convTransposeB_CP_4758_elements(43), ack => convTransposeB_CP_4758_elements(83), clk => clk, reset =>reset);
    -- CP-element group 84:  transition  output  delay-element  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	43 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (4) 
      -- CP-element group 84: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1969/$exit
      -- CP-element group 84: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1973_konst_delay_trans
      -- CP-element group 84: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_req
      -- 
    phi_stmt_1969_req_5488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1969_req_5488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(84), ack => phi_stmt_1969_req_0); -- 
    -- Element group convTransposeB_CP_4758_elements(84) is a control-delay.
    cp_element_84_delay: control_delay_element  generic map(name => " 84_delay", delay_value => 1)  port map(req => convTransposeB_CP_4758_elements(43), ack => convTransposeB_CP_4758_elements(84), clk => clk, reset =>reset);
    -- CP-element group 85:  join  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	81 
    -- CP-element group 85: 	82 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	99 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1854/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(81) & convTransposeB_CP_4758_elements(82) & convTransposeB_CP_4758_elements(83) & convTransposeB_CP_4758_elements(84);
      gj_convTransposeB_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1995/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1995/SplitProtocol/Sample/ra
      -- 
    ra_5508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1995_inst_ack_0, ack => convTransposeB_CP_4758_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1995/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1995/SplitProtocol/Update/ca
      -- 
    ca_5513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1995_inst_ack_1, ack => convTransposeB_CP_4758_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	98 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1990/$exit
      -- CP-element group 88: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1995/$exit
      -- CP-element group 88: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1995/SplitProtocol/$exit
      -- CP-element group 88: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1990/phi_stmt_1990_req
      -- 
    phi_stmt_1990_req_5514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1990_req_5514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(88), ack => phi_stmt_1990_req_1); -- 
    convTransposeB_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(86) & convTransposeB_CP_4758_elements(87);
      gj_convTransposeB_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/SplitProtocol/Sample/ra
      -- 
    ra_5531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1986_inst_ack_0, ack => convTransposeB_CP_4758_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/SplitProtocol/Update/ca
      -- 
    ca_5536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1986_inst_ack_1, ack => convTransposeB_CP_4758_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	98 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/$exit
      -- CP-element group 91: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/$exit
      -- CP-element group 91: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_req
      -- 
    phi_stmt_1983_req_5537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1983_req_5537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(91), ack => phi_stmt_1983_req_0); -- 
    convTransposeB_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(89) & convTransposeB_CP_4758_elements(90);
      gj_convTransposeB_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/SplitProtocol/Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/SplitProtocol/Sample/ra
      -- 
    ra_5554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1982_inst_ack_0, ack => convTransposeB_CP_4758_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/SplitProtocol/Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/SplitProtocol/Update/ca
      -- 
    ca_5559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1982_inst_ack_1, ack => convTransposeB_CP_4758_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	98 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/$exit
      -- CP-element group 94: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/$exit
      -- CP-element group 94: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/SplitProtocol/$exit
      -- CP-element group 94: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_req
      -- 
    phi_stmt_1976_req_5560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1976_req_5560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(94), ack => phi_stmt_1976_req_1); -- 
    convTransposeB_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(92) & convTransposeB_CP_4758_elements(93);
      gj_convTransposeB_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/SplitProtocol/Sample/ra
      -- 
    ra_5577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1975_inst_ack_0, ack => convTransposeB_CP_4758_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/SplitProtocol/Update/ca
      -- 
    ca_5582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1975_inst_ack_1, ack => convTransposeB_CP_4758_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/$exit
      -- CP-element group 97: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/$exit
      -- CP-element group 97: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_req
      -- 
    phi_stmt_1969_req_5583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1969_req_5583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(97), ack => phi_stmt_1969_req_1); -- 
    convTransposeB_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(95) & convTransposeB_CP_4758_elements(96);
      gj_convTransposeB_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	88 
    -- CP-element group 98: 	91 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1854/ifx_xend128_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(88) & convTransposeB_CP_4758_elements(91) & convTransposeB_CP_4758_elements(94) & convTransposeB_CP_4758_elements(97);
      gj_convTransposeB_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  merge  fork  transition  place  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	85 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	101 
    -- CP-element group 99: 	102 
    -- CP-element group 99: 	103 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1854/merge_stmt_1968_PhiReqMerge
      -- CP-element group 99: 	 branch_block_stmt_1854/merge_stmt_1968_PhiAck/$entry
      -- 
    convTransposeB_CP_4758_elements(99) <= OrReduce(convTransposeB_CP_4758_elements(85) & convTransposeB_CP_4758_elements(98));
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1854/merge_stmt_1968_PhiAck/phi_stmt_1969_ack
      -- 
    phi_stmt_1969_ack_5588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1969_ack_0, ack => convTransposeB_CP_4758_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1854/merge_stmt_1968_PhiAck/phi_stmt_1976_ack
      -- 
    phi_stmt_1976_ack_5589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1976_ack_0, ack => convTransposeB_CP_4758_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_1854/merge_stmt_1968_PhiAck/phi_stmt_1983_ack
      -- 
    phi_stmt_1983_ack_5590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1983_ack_0, ack => convTransposeB_CP_4758_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	99 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1854/merge_stmt_1968_PhiAck/phi_stmt_1990_ack
      -- 
    phi_stmt_1990_ack_5591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1990_ack_0, ack => convTransposeB_CP_4758_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  place  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	101 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	44 
    -- CP-element group 104: 	45 
    -- CP-element group 104: 	46 
    -- CP-element group 104: 	47 
    -- CP-element group 104: 	48 
    -- CP-element group 104: 	49 
    -- CP-element group 104: 	50 
    -- CP-element group 104: 	51 
    -- CP-element group 104: 	53 
    -- CP-element group 104: 	55 
    -- CP-element group 104: 	57 
    -- CP-element group 104: 	60 
    -- CP-element group 104: 	62 
    -- CP-element group 104: 	65 
    -- CP-element group 104: 	66 
    -- CP-element group 104: 	67 
    -- CP-element group 104:  members (56) 
      -- CP-element group 104: 	 branch_block_stmt_1854/merge_stmt_1968__exit__
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118__entry__
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2030_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2030_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/$entry
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2030_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2030_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2030_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2030_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2034_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2034_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2034_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2034_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2034_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2034_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2038_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2038_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2038_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2038_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2038_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2038_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2068_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2068_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2068_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2068_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2068_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2068_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2075_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2074_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2075_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2075_complete/req
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2079_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2098_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/array_obj_ref_2097_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2098_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/addr_of_2098_complete/req
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/ptr_deref_2101_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2106_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2106_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2106_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2106_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2106_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1854/assign_stmt_2002_to_assign_stmt_2118/type_cast_2106_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1854/merge_stmt_1968_PhiAck/$exit
      -- 
    rr_5092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => type_cast_2030_inst_req_0); -- 
    cr_5097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => type_cast_2030_inst_req_1); -- 
    rr_5106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => type_cast_2034_inst_req_0); -- 
    cr_5111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => type_cast_2034_inst_req_1); -- 
    rr_5120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => type_cast_2038_inst_req_0); -- 
    cr_5125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => type_cast_2038_inst_req_1); -- 
    rr_5134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => type_cast_2068_inst_req_0); -- 
    cr_5139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => type_cast_2068_inst_req_1); -- 
    req_5170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => array_obj_ref_2074_index_offset_req_1); -- 
    req_5185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => addr_of_2075_final_reg_req_1); -- 
    cr_5230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => ptr_deref_2079_load_0_req_1); -- 
    req_5266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => array_obj_ref_2097_index_offset_req_1); -- 
    req_5281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => addr_of_2098_final_reg_req_1); -- 
    cr_5331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => ptr_deref_2101_store_0_req_1); -- 
    rr_5340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => type_cast_2106_inst_req_0); -- 
    cr_5345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => type_cast_2106_inst_req_1); -- 
    convTransposeB_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(100) & convTransposeB_CP_4758_elements(101) & convTransposeB_CP_4758_elements(102) & convTransposeB_CP_4758_elements(103);
      gj_convTransposeB_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	76 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2195/SplitProtocol/Sample/ra
      -- CP-element group 105: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2195/SplitProtocol/Sample/$exit
      -- 
    ra_5635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2195_inst_ack_0, ack => convTransposeB_CP_4758_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2195/SplitProtocol/Update/ca
      -- CP-element group 106: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2195/SplitProtocol/Update/$exit
      -- 
    ca_5640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2195_inst_ack_1, ack => convTransposeB_CP_4758_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	112 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2190/$exit
      -- CP-element group 107: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_req
      -- CP-element group 107: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2195/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2195/$exit
      -- 
    phi_stmt_2190_req_5641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2190_req_5641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(107), ack => phi_stmt_2190_req_1); -- 
    convTransposeB_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(105) & convTransposeB_CP_4758_elements(106);
      gj_convTransposeB_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  transition  output  delay-element  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	76 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	112 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_req
      -- CP-element group 108: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2183_konst_delay_trans
      -- CP-element group 108: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/$exit
      -- 
    phi_stmt_2177_req_5649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2177_req_5649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(108), ack => phi_stmt_2177_req_1); -- 
    -- Element group convTransposeB_CP_4758_elements(108) is a control-delay.
    cp_element_108_delay: control_delay_element  generic map(name => " 108_delay", delay_value => 1)  port map(req => convTransposeB_CP_4758_elements(76), ack => convTransposeB_CP_4758_elements(108), clk => clk, reset =>reset);
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/SplitProtocol/Sample/ra
      -- CP-element group 109: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/SplitProtocol/Sample/$exit
      -- 
    ra_5666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2189_inst_ack_0, ack => convTransposeB_CP_4758_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	76 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/SplitProtocol/Update/ca
      -- 
    ca_5671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2189_inst_ack_1, ack => convTransposeB_CP_4758_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/$exit
      -- CP-element group 111: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/$exit
      -- CP-element group 111: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_req
      -- 
    phi_stmt_2184_req_5672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2184_req_5672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(111), ack => phi_stmt_2184_req_1); -- 
    convTransposeB_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(109) & convTransposeB_CP_4758_elements(110);
      gj_convTransposeB_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	107 
    -- CP-element group 112: 	108 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	123 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_1854/ifx_xelse_ifx_xend128_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(107) & convTransposeB_CP_4758_elements(108) & convTransposeB_CP_4758_elements(111);
      gj_convTransposeB_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	69 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Sample/ra
      -- CP-element group 113: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Sample/$exit
      -- 
    ra_5692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2193_inst_ack_0, ack => convTransposeB_CP_4758_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Update/ca
      -- 
    ca_5697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2193_inst_ack_1, ack => convTransposeB_CP_4758_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	122 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/$exit
      -- CP-element group 115: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/$exit
      -- CP-element group 115: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2190/$exit
      -- CP-element group 115: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2190/phi_stmt_2190_req
      -- 
    phi_stmt_2190_req_5698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2190_req_5698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(115), ack => phi_stmt_2190_req_0); -- 
    convTransposeB_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(113) & convTransposeB_CP_4758_elements(114);
      gj_convTransposeB_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Sample/ra
      -- CP-element group 116: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Sample/$exit
      -- 
    ra_5715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2180_inst_ack_0, ack => convTransposeB_CP_4758_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Update/ca
      -- CP-element group 117: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Update/$exit
      -- 
    ca_5720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2180_inst_ack_1, ack => convTransposeB_CP_4758_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	122 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_req
      -- CP-element group 118: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/$exit
      -- CP-element group 118: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/$exit
      -- 
    phi_stmt_2177_req_5721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2177_req_5721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(118), ack => phi_stmt_2177_req_0); -- 
    convTransposeB_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(116) & convTransposeB_CP_4758_elements(117);
      gj_convTransposeB_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	69 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/SplitProtocol/Sample/ra
      -- CP-element group 119: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/SplitProtocol/Sample/$exit
      -- 
    ra_5738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2187_inst_ack_0, ack => convTransposeB_CP_4758_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	69 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/SplitProtocol/Update/ca
      -- CP-element group 120: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/SplitProtocol/Update/$exit
      -- 
    ca_5743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2187_inst_ack_1, ack => convTransposeB_CP_4758_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_req
      -- CP-element group 121: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/$exit
      -- CP-element group 121: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/$exit
      -- CP-element group 121: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/$exit
      -- 
    phi_stmt_2184_req_5744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2184_req_5744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(121), ack => phi_stmt_2184_req_0); -- 
    convTransposeB_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(119) & convTransposeB_CP_4758_elements(120);
      gj_convTransposeB_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	115 
    -- CP-element group 122: 	118 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1854/ifx_xthen_ifx_xend128_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(115) & convTransposeB_CP_4758_elements(118) & convTransposeB_CP_4758_elements(121);
      gj_convTransposeB_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  fork  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	112 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	126 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1854/merge_stmt_2176_PhiAck/$entry
      -- CP-element group 123: 	 branch_block_stmt_1854/merge_stmt_2176_PhiReqMerge
      -- 
    convTransposeB_CP_4758_elements(123) <= OrReduce(convTransposeB_CP_4758_elements(112) & convTransposeB_CP_4758_elements(122));
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	127 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1854/merge_stmt_2176_PhiAck/phi_stmt_2177_ack
      -- 
    phi_stmt_2177_ack_5749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2177_ack_0, ack => convTransposeB_CP_4758_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1854/merge_stmt_2176_PhiAck/phi_stmt_2184_ack
      -- 
    phi_stmt_2184_ack_5750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2184_ack_0, ack => convTransposeB_CP_4758_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	123 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_1854/merge_stmt_2176_PhiAck/phi_stmt_2190_ack
      -- 
    phi_stmt_2190_ack_5751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2190_ack_0, ack => convTransposeB_CP_4758_elements(126)); -- 
    -- CP-element group 127:  join  transition  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	124 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_1854/merge_stmt_2176_PhiAck/$exit
      -- 
    convTransposeB_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(124) & convTransposeB_CP_4758_elements(125) & convTransposeB_CP_4758_elements(126);
      gj_convTransposeB_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(127), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom86_2096_resized : std_logic_vector(13 downto 0);
    signal R_idxprom86_2096_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2073_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2073_scaled : std_logic_vector(13 downto 0);
    signal add45_1928 : std_logic_vector(15 downto 0);
    signal add58_1939 : std_logic_vector(15 downto 0);
    signal add77_2049 : std_logic_vector(63 downto 0);
    signal add79_2059 : std_logic_vector(63 downto 0);
    signal add91_2113 : std_logic_vector(31 downto 0);
    signal add98_2131 : std_logic_vector(15 downto 0);
    signal add_1906 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2007 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2074_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2074_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2074_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2074_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2074_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2074_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2097_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2097_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2097_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2097_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2097_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2097_root_address : std_logic_vector(13 downto 0);
    signal arrayidx82_2076 : std_logic_vector(31 downto 0);
    signal arrayidx87_2099 : std_logic_vector(31 downto 0);
    signal call11_1875 : std_logic_vector(15 downto 0);
    signal call13_1878 : std_logic_vector(15 downto 0);
    signal call14_1881 : std_logic_vector(15 downto 0);
    signal call15_1884 : std_logic_vector(15 downto 0);
    signal call16_1897 : std_logic_vector(15 downto 0);
    signal call18_1909 : std_logic_vector(15 downto 0);
    signal call1_1860 : std_logic_vector(15 downto 0);
    signal call20_1912 : std_logic_vector(15 downto 0);
    signal call22_1915 : std_logic_vector(15 downto 0);
    signal call3_1863 : std_logic_vector(15 downto 0);
    signal call5_1866 : std_logic_vector(15 downto 0);
    signal call7_1869 : std_logic_vector(15 downto 0);
    signal call9_1872 : std_logic_vector(15 downto 0);
    signal call_1857 : std_logic_vector(15 downto 0);
    signal cmp106_2144 : std_logic_vector(0 downto 0);
    signal cmp117_2169 : std_logic_vector(0 downto 0);
    signal cmp_2118 : std_logic_vector(0 downto 0);
    signal conv112_2164 : std_logic_vector(31 downto 0);
    signal conv115_1960 : std_logic_vector(31 downto 0);
    signal conv17_1901 : std_logic_vector(31 downto 0);
    signal conv65_2031 : std_logic_vector(63 downto 0);
    signal conv68_1948 : std_logic_vector(63 downto 0);
    signal conv70_2035 : std_logic_vector(63 downto 0);
    signal conv73_1952 : std_logic_vector(63 downto 0);
    signal conv75_2039 : std_logic_vector(63 downto 0);
    signal conv90_2107 : std_logic_vector(31 downto 0);
    signal conv94_1956 : std_logic_vector(31 downto 0);
    signal conv_1888 : std_logic_vector(31 downto 0);
    signal idxprom86_2092 : std_logic_vector(63 downto 0);
    signal idxprom_2069 : std_logic_vector(63 downto 0);
    signal inc110_2148 : std_logic_vector(15 downto 0);
    signal inc110x_xinput_dim0x_x2_2153 : std_logic_vector(15 downto 0);
    signal inc_2139 : std_logic_vector(15 downto 0);
    signal indvar_1969 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2202 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2190 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1990 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2184 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1983 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2160 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2177 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1976 : std_logic_vector(15 downto 0);
    signal mul54_2022 : std_logic_vector(15 downto 0);
    signal mul76_2044 : std_logic_vector(63 downto 0);
    signal mul78_2054 : std_logic_vector(63 downto 0);
    signal mul_2012 : std_logic_vector(15 downto 0);
    signal ptr_deref_2079_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2079_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2079_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2079_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2079_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2101_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2101_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2101_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2101_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2101_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2101_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1894 : std_logic_vector(31 downto 0);
    signal shr116132_1966 : std_logic_vector(31 downto 0);
    signal shr131_1922 : std_logic_vector(15 downto 0);
    signal shr81_2065 : std_logic_vector(31 downto 0);
    signal shr85_2086 : std_logic_vector(63 downto 0);
    signal sub48_2017 : std_logic_vector(15 downto 0);
    signal sub61_1944 : std_logic_vector(15 downto 0);
    signal sub62_2027 : std_logic_vector(15 downto 0);
    signal sub_1933 : std_logic_vector(15 downto 0);
    signal tmp1_2002 : std_logic_vector(31 downto 0);
    signal tmp83_2080 : std_logic_vector(63 downto 0);
    signal type_cast_1892_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1920_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1926_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1937_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1964_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1973_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1975_wire : std_logic_vector(31 downto 0);
    signal type_cast_1980_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1982_wire : std_logic_vector(15 downto 0);
    signal type_cast_1986_wire : std_logic_vector(15 downto 0);
    signal type_cast_1989_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1993_wire : std_logic_vector(15 downto 0);
    signal type_cast_1995_wire : std_logic_vector(15 downto 0);
    signal type_cast_2000_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2063_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2084_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2090_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2111_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2129_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2137_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2157_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2180_wire : std_logic_vector(15 downto 0);
    signal type_cast_2183_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2187_wire : std_logic_vector(15 downto 0);
    signal type_cast_2189_wire : std_logic_vector(15 downto 0);
    signal type_cast_2193_wire : std_logic_vector(15 downto 0);
    signal type_cast_2195_wire : std_logic_vector(15 downto 0);
    signal type_cast_2200_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2208_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2074_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2074_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2074_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2074_resized_base_address <= "00000000000000";
    array_obj_ref_2097_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2097_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2097_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2097_resized_base_address <= "00000000000000";
    ptr_deref_2079_word_offset_0 <= "00000000000000";
    ptr_deref_2101_word_offset_0 <= "00000000000000";
    type_cast_1892_wire_constant <= "00000000000000000000000000010000";
    type_cast_1920_wire_constant <= "0000000000000010";
    type_cast_1926_wire_constant <= "1111111111111111";
    type_cast_1937_wire_constant <= "1111111111111111";
    type_cast_1964_wire_constant <= "00000000000000000000000000000001";
    type_cast_1973_wire_constant <= "00000000000000000000000000000000";
    type_cast_1980_wire_constant <= "0000000000000000";
    type_cast_1989_wire_constant <= "0000000000000000";
    type_cast_2000_wire_constant <= "00000000000000000000000000000100";
    type_cast_2063_wire_constant <= "00000000000000000000000000000010";
    type_cast_2084_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2090_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2111_wire_constant <= "00000000000000000000000000000100";
    type_cast_2129_wire_constant <= "0000000000000100";
    type_cast_2137_wire_constant <= "0000000000000001";
    type_cast_2157_wire_constant <= "0000000000000000";
    type_cast_2183_wire_constant <= "0000000000000000";
    type_cast_2200_wire_constant <= "00000000000000000000000000000001";
    type_cast_2208_wire_constant <= "0000000000000001";
    phi_stmt_1969: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1973_wire_constant & type_cast_1975_wire;
      req <= phi_stmt_1969_req_0 & phi_stmt_1969_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1969",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1969_ack_0,
          idata => idata,
          odata => indvar_1969,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1969
    phi_stmt_1976: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1980_wire_constant & type_cast_1982_wire;
      req <= phi_stmt_1976_req_0 & phi_stmt_1976_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1976",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1976_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1976,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1976
    phi_stmt_1983: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1986_wire & type_cast_1989_wire_constant;
      req <= phi_stmt_1983_req_0 & phi_stmt_1983_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1983",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1983_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1983,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1983
    phi_stmt_1990: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1993_wire & type_cast_1995_wire;
      req <= phi_stmt_1990_req_0 & phi_stmt_1990_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1990",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1990_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1990,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1990
    phi_stmt_2177: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2180_wire & type_cast_2183_wire_constant;
      req <= phi_stmt_2177_req_0 & phi_stmt_2177_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2177",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2177_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2177,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2177
    phi_stmt_2184: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2187_wire & type_cast_2189_wire;
      req <= phi_stmt_2184_req_0 & phi_stmt_2184_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2184",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2184_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2184,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2184
    phi_stmt_2190: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2193_wire & type_cast_2195_wire;
      req <= phi_stmt_2190_req_0 & phi_stmt_2190_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2190",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2190_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2190,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2190
    -- flow-through select operator MUX_2159_inst
    input_dim1x_x2_2160 <= type_cast_2157_wire_constant when (cmp106_2144(0) /=  '0') else inc_2139;
    addr_of_2075_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2075_final_reg_req_0;
      addr_of_2075_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2075_final_reg_req_1;
      addr_of_2075_final_reg_ack_1<= rack(0);
      addr_of_2075_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2075_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2074_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_2076,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2098_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2098_final_reg_req_0;
      addr_of_2098_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2098_final_reg_req_1;
      addr_of_2098_final_reg_ack_1<= rack(0);
      addr_of_2098_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2098_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2097_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2099,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1887_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1887_inst_req_0;
      type_cast_1887_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1887_inst_req_1;
      type_cast_1887_inst_ack_1<= rack(0);
      type_cast_1887_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1887_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1884,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1888,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1900_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1900_inst_req_0;
      type_cast_1900_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1900_inst_req_1;
      type_cast_1900_inst_ack_1<= rack(0);
      type_cast_1900_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1900_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1897,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1901,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1947_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1947_inst_req_0;
      type_cast_1947_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1947_inst_req_1;
      type_cast_1947_inst_ack_1<= rack(0);
      type_cast_1947_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1947_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1915,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_1948,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1951_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1951_inst_req_0;
      type_cast_1951_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1951_inst_req_1;
      type_cast_1951_inst_ack_1<= rack(0);
      type_cast_1951_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1951_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1912,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_1952,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1955_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1955_inst_req_0;
      type_cast_1955_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1955_inst_req_1;
      type_cast_1955_inst_ack_1<= rack(0);
      type_cast_1955_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1955_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1863,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_1956,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1959_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1959_inst_req_0;
      type_cast_1959_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1959_inst_req_1;
      type_cast_1959_inst_ack_1<= rack(0);
      type_cast_1959_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1959_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1857,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_1960,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1975_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1975_inst_req_0;
      type_cast_1975_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1975_inst_req_1;
      type_cast_1975_inst_ack_1<= rack(0);
      type_cast_1975_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1975_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2202,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1975_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1982_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1982_inst_req_0;
      type_cast_1982_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1982_inst_req_1;
      type_cast_1982_inst_ack_1<= rack(0);
      type_cast_1982_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1982_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2177,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1982_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1986_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1986_inst_req_0;
      type_cast_1986_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1986_inst_req_1;
      type_cast_1986_inst_ack_1<= rack(0);
      type_cast_1986_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1986_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2184,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1986_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1993_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1993_inst_req_0;
      type_cast_1993_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1993_inst_req_1;
      type_cast_1993_inst_ack_1<= rack(0);
      type_cast_1993_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1993_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr131_1922,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1993_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1995_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1995_inst_req_0;
      type_cast_1995_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1995_inst_req_1;
      type_cast_1995_inst_ack_1<= rack(0);
      type_cast_1995_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1995_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2190,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1995_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2030_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2030_inst_req_0;
      type_cast_2030_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2030_inst_req_1;
      type_cast_2030_inst_ack_1<= rack(0);
      type_cast_2030_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2030_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1976,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2031,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2034_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2034_inst_req_0;
      type_cast_2034_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2034_inst_req_1;
      type_cast_2034_inst_ack_1<= rack(0);
      type_cast_2034_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2034_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub62_2027,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2035,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2038_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2038_inst_req_0;
      type_cast_2038_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2038_inst_req_1;
      type_cast_2038_inst_ack_1<= rack(0);
      type_cast_2038_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2038_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub48_2017,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2039,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2068_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2068_inst_req_0;
      type_cast_2068_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2068_inst_req_1;
      type_cast_2068_inst_ack_1<= rack(0);
      type_cast_2068_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2068_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr81_2065,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2069,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2106_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2106_inst_req_0;
      type_cast_2106_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2106_inst_req_1;
      type_cast_2106_inst_ack_1<= rack(0);
      type_cast_2106_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2106_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1976,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_2107,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2147_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2147_inst_req_0;
      type_cast_2147_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2147_inst_req_1;
      type_cast_2147_inst_ack_1<= rack(0);
      type_cast_2147_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2147_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp106_2144,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc110_2148,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2163_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2163_inst_req_0;
      type_cast_2163_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2163_inst_req_1;
      type_cast_2163_inst_ack_1<= rack(0);
      type_cast_2163_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2163_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2153,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_2164,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2180_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2180_inst_req_0;
      type_cast_2180_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2180_inst_req_1;
      type_cast_2180_inst_ack_1<= rack(0);
      type_cast_2180_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2180_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add98_2131,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2180_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2187_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2187_inst_req_0;
      type_cast_2187_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2187_inst_req_1;
      type_cast_2187_inst_ack_1<= rack(0);
      type_cast_2187_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2187_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1983,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2187_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2189_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2189_inst_req_0;
      type_cast_2189_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2189_inst_req_1;
      type_cast_2189_inst_ack_1<= rack(0);
      type_cast_2189_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2189_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2160,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2189_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2193_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2193_inst_req_0;
      type_cast_2193_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2193_inst_req_1;
      type_cast_2193_inst_ack_1<= rack(0);
      type_cast_2193_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2193_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1990,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2193_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2195_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2195_inst_req_0;
      type_cast_2195_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2195_inst_req_1;
      type_cast_2195_inst_ack_1<= rack(0);
      type_cast_2195_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2195_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2153,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2195_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2074_index_1_rename
    process(R_idxprom_2073_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2073_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2073_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2074_index_1_resize
    process(idxprom_2069) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2069;
      ov := iv(13 downto 0);
      R_idxprom_2073_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2074_root_address_inst
    process(array_obj_ref_2074_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2074_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2074_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2097_index_1_rename
    process(R_idxprom86_2096_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom86_2096_resized;
      ov(13 downto 0) := iv;
      R_idxprom86_2096_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2097_index_1_resize
    process(idxprom86_2092) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom86_2092;
      ov := iv(13 downto 0);
      R_idxprom86_2096_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2097_root_address_inst
    process(array_obj_ref_2097_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2097_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2097_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2079_addr_0
    process(ptr_deref_2079_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2079_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2079_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2079_base_resize
    process(arrayidx82_2076) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_2076;
      ov := iv(13 downto 0);
      ptr_deref_2079_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2079_gather_scatter
    process(ptr_deref_2079_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2079_data_0;
      ov(63 downto 0) := iv;
      tmp83_2080 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2079_root_address_inst
    process(ptr_deref_2079_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2079_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2079_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2101_addr_0
    process(ptr_deref_2101_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2101_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2101_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2101_base_resize
    process(arrayidx87_2099) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2099;
      ov := iv(13 downto 0);
      ptr_deref_2101_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2101_gather_scatter
    process(tmp83_2080) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp83_2080;
      ov(63 downto 0) := iv;
      ptr_deref_2101_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2101_root_address_inst
    process(ptr_deref_2101_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2101_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2101_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2119_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2118;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2119_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2119_branch_req_0,
          ack0 => if_stmt_2119_branch_ack_0,
          ack1 => if_stmt_2119_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2170_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp117_2169;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2170_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2170_branch_req_0,
          ack0 => if_stmt_2170_branch_ack_0,
          ack1 => if_stmt_2170_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1927_inst
    process(call7_1869) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1869, type_cast_1926_wire_constant, tmp_var);
      add45_1928 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1938_inst
    process(call9_1872) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1872, type_cast_1937_wire_constant, tmp_var);
      add58_1939 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2016_inst
    process(sub_1933, mul_2012) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1933, mul_2012, tmp_var);
      sub48_2017 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2026_inst
    process(sub61_1944, mul54_2022) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub61_1944, mul54_2022, tmp_var);
      sub62_2027 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2130_inst
    process(input_dim2x_x1_1976) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1976, type_cast_2129_wire_constant, tmp_var);
      add98_2131 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2138_inst
    process(input_dim1x_x1_1983) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1983, type_cast_2137_wire_constant, tmp_var);
      inc_2139 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2152_inst
    process(inc110_2148, input_dim0x_x2_1990) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc110_2148, input_dim0x_x2_1990, tmp_var);
      inc110x_xinput_dim0x_x2_2153 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2006_inst
    process(add_1906, tmp1_2002) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1906, tmp1_2002, tmp_var);
      add_src_0x_x0_2007 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2112_inst
    process(conv90_2107) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv90_2107, type_cast_2111_wire_constant, tmp_var);
      add91_2113 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2201_inst
    process(indvar_1969) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1969, type_cast_2200_wire_constant, tmp_var);
      indvarx_xnext_2202 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2048_inst
    process(mul76_2044, conv70_2035) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul76_2044, conv70_2035, tmp_var);
      add77_2049 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2058_inst
    process(mul78_2054, conv65_2031) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul78_2054, conv65_2031, tmp_var);
      add79_2059 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2091_inst
    process(shr85_2086) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr85_2086, type_cast_2090_wire_constant, tmp_var);
      idxprom86_2092 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2143_inst
    process(inc_2139, call1_1860) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2139, call1_1860, tmp_var);
      cmp106_2144 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2168_inst
    process(conv112_2164, shr116132_1966) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv112_2164, shr116132_1966, tmp_var);
      cmp117_2169 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1921_inst
    process(call_1857) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1857, type_cast_1920_wire_constant, tmp_var);
      shr131_1922 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1965_inst
    process(conv115_1960) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_1960, type_cast_1964_wire_constant, tmp_var);
      shr116132_1966 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2064_inst
    process(add_src_0x_x0_2007) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2007, type_cast_2063_wire_constant, tmp_var);
      shr81_2065 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2085_inst
    process(add79_2059) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_2059, type_cast_2084_wire_constant, tmp_var);
      shr85_2086 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2011_inst
    process(input_dim0x_x2_1990, call13_1878) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_1990, call13_1878, tmp_var);
      mul_2012 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2021_inst
    process(input_dim1x_x1_1983, call13_1878) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1983, call13_1878, tmp_var);
      mul54_2022 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2001_inst
    process(indvar_1969) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1969, type_cast_2000_wire_constant, tmp_var);
      tmp1_2002 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2043_inst
    process(conv75_2039, conv73_1952) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv75_2039, conv73_1952, tmp_var);
      mul76_2044 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2053_inst
    process(add77_2049, conv68_1948) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add77_2049, conv68_1948, tmp_var);
      mul78_2054 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1905_inst
    process(shl_1894, conv17_1901) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1894, conv17_1901, tmp_var);
      add_1906 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1893_inst
    process(conv_1888) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1888, type_cast_1892_wire_constant, tmp_var);
      shl_1894 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1932_inst
    process(add45_1928, call14_1881) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add45_1928, call14_1881, tmp_var);
      sub_1933 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1943_inst
    process(add58_1939, call14_1881) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add58_1939, call14_1881, tmp_var);
      sub61_1944 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2117_inst
    process(add91_2113, conv94_1956) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add91_2113, conv94_1956, tmp_var);
      cmp_2118 <= tmp_var; --
    end process;
    -- shared split operator group (29) : array_obj_ref_2074_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2073_scaled;
      array_obj_ref_2074_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2074_index_offset_req_0;
      array_obj_ref_2074_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2074_index_offset_req_1;
      array_obj_ref_2074_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : array_obj_ref_2097_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom86_2096_scaled;
      array_obj_ref_2097_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2097_index_offset_req_0;
      array_obj_ref_2097_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2097_index_offset_req_1;
      array_obj_ref_2097_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared load operator group (0) : ptr_deref_2079_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2079_load_0_req_0;
      ptr_deref_2079_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2079_load_0_req_1;
      ptr_deref_2079_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2079_word_address_0;
      ptr_deref_2079_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2101_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2101_store_0_req_0;
      ptr_deref_2101_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2101_store_0_req_1;
      ptr_deref_2101_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2101_word_address_0;
      data_in <= ptr_deref_2101_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1914_inst RPIPE_Block1_start_1911_inst RPIPE_Block1_start_1908_inst RPIPE_Block1_start_1896_inst RPIPE_Block1_start_1883_inst RPIPE_Block1_start_1880_inst RPIPE_Block1_start_1877_inst RPIPE_Block1_start_1874_inst RPIPE_Block1_start_1871_inst RPIPE_Block1_start_1868_inst RPIPE_Block1_start_1865_inst RPIPE_Block1_start_1862_inst RPIPE_Block1_start_1859_inst RPIPE_Block1_start_1856_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block1_start_1914_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block1_start_1911_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block1_start_1908_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block1_start_1896_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block1_start_1883_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block1_start_1880_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block1_start_1877_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block1_start_1874_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block1_start_1871_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block1_start_1868_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block1_start_1865_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block1_start_1862_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block1_start_1859_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block1_start_1856_inst_req_0;
      RPIPE_Block1_start_1914_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block1_start_1911_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block1_start_1908_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block1_start_1896_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block1_start_1883_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block1_start_1880_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block1_start_1877_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block1_start_1874_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block1_start_1871_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block1_start_1868_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block1_start_1865_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block1_start_1862_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block1_start_1859_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block1_start_1856_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block1_start_1914_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block1_start_1911_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block1_start_1908_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block1_start_1896_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block1_start_1883_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block1_start_1880_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block1_start_1877_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block1_start_1874_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block1_start_1871_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block1_start_1868_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block1_start_1865_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block1_start_1862_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block1_start_1859_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block1_start_1856_inst_req_1;
      RPIPE_Block1_start_1914_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block1_start_1911_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block1_start_1908_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block1_start_1896_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block1_start_1883_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block1_start_1880_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block1_start_1877_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block1_start_1874_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block1_start_1871_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block1_start_1868_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block1_start_1865_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block1_start_1862_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block1_start_1859_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block1_start_1856_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call22_1915 <= data_out(223 downto 208);
      call20_1912 <= data_out(207 downto 192);
      call18_1909 <= data_out(191 downto 176);
      call16_1897 <= data_out(175 downto 160);
      call15_1884 <= data_out(159 downto 144);
      call14_1881 <= data_out(143 downto 128);
      call13_1878 <= data_out(127 downto 112);
      call11_1875 <= data_out(111 downto 96);
      call9_1872 <= data_out(95 downto 80);
      call7_1869 <= data_out(79 downto 64);
      call5_1866 <= data_out(63 downto 48);
      call3_1863 <= data_out(47 downto 32);
      call1_1860 <= data_out(31 downto 16);
      call_1857 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_2206_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_2206_inst_req_0;
      WPIPE_Block1_done_2206_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_2206_inst_req_1;
      WPIPE_Block1_done_2206_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2208_wire_constant;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_5768_start: Boolean;
  signal convTransposeC_CP_5768_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block2_start_2226_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2229_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2241_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2226_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2275_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2238_inst_ack_1 : boolean;
  signal type_cast_2248_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2241_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2269_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2275_inst_ack_0 : boolean;
  signal type_cast_2248_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2269_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2244_inst_req_0 : boolean;
  signal type_cast_2312_inst_ack_0 : boolean;
  signal type_cast_2248_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2244_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2229_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2235_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2244_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2232_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2235_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2241_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2238_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2238_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2235_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2257_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2257_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2272_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2235_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2241_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2244_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2232_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2229_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2232_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2226_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2257_inst_req_1 : boolean;
  signal type_cast_2261_inst_ack_1 : boolean;
  signal type_cast_2261_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2269_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2257_inst_ack_1 : boolean;
  signal type_cast_2248_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2269_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2232_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2275_inst_req_1 : boolean;
  signal type_cast_2261_inst_req_1 : boolean;
  signal type_cast_2261_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2272_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2275_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2226_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2272_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2238_inst_req_1 : boolean;
  signal type_cast_2402_inst_ack_0 : boolean;
  signal type_cast_2402_inst_req_1 : boolean;
  signal type_cast_2320_inst_req_1 : boolean;
  signal type_cast_2320_inst_ack_1 : boolean;
  signal type_cast_2308_inst_ack_1 : boolean;
  signal type_cast_2320_inst_req_0 : boolean;
  signal type_cast_2320_inst_ack_0 : boolean;
  signal type_cast_2308_inst_req_1 : boolean;
  signal type_cast_2312_inst_ack_1 : boolean;
  signal type_cast_2316_inst_req_1 : boolean;
  signal type_cast_2316_inst_ack_1 : boolean;
  signal type_cast_2312_inst_req_1 : boolean;
  signal type_cast_2402_inst_req_0 : boolean;
  signal type_cast_2308_inst_ack_0 : boolean;
  signal type_cast_2308_inst_req_0 : boolean;
  signal type_cast_2316_inst_req_0 : boolean;
  signal type_cast_2316_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2272_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2229_inst_req_0 : boolean;
  signal type_cast_2312_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2223_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2223_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2217_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2217_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2217_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2217_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2220_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2220_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2220_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2220_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2223_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2223_inst_ack_0 : boolean;
  signal type_cast_2402_inst_ack_1 : boolean;
  signal type_cast_2406_inst_req_0 : boolean;
  signal type_cast_2406_inst_ack_0 : boolean;
  signal type_cast_2406_inst_req_1 : boolean;
  signal type_cast_2406_inst_ack_1 : boolean;
  signal type_cast_2410_inst_req_0 : boolean;
  signal type_cast_2410_inst_ack_0 : boolean;
  signal type_cast_2410_inst_req_1 : boolean;
  signal type_cast_2410_inst_ack_1 : boolean;
  signal type_cast_2440_inst_req_0 : boolean;
  signal type_cast_2440_inst_ack_0 : boolean;
  signal type_cast_2440_inst_req_1 : boolean;
  signal type_cast_2440_inst_ack_1 : boolean;
  signal array_obj_ref_2446_index_offset_req_0 : boolean;
  signal array_obj_ref_2446_index_offset_ack_0 : boolean;
  signal array_obj_ref_2446_index_offset_req_1 : boolean;
  signal array_obj_ref_2446_index_offset_ack_1 : boolean;
  signal addr_of_2447_final_reg_req_0 : boolean;
  signal addr_of_2447_final_reg_ack_0 : boolean;
  signal addr_of_2447_final_reg_req_1 : boolean;
  signal addr_of_2447_final_reg_ack_1 : boolean;
  signal ptr_deref_2451_load_0_req_0 : boolean;
  signal ptr_deref_2451_load_0_ack_0 : boolean;
  signal ptr_deref_2451_load_0_req_1 : boolean;
  signal ptr_deref_2451_load_0_ack_1 : boolean;
  signal array_obj_ref_2469_index_offset_req_0 : boolean;
  signal array_obj_ref_2469_index_offset_ack_0 : boolean;
  signal array_obj_ref_2469_index_offset_req_1 : boolean;
  signal array_obj_ref_2469_index_offset_ack_1 : boolean;
  signal addr_of_2470_final_reg_req_0 : boolean;
  signal addr_of_2470_final_reg_ack_0 : boolean;
  signal addr_of_2470_final_reg_req_1 : boolean;
  signal addr_of_2470_final_reg_ack_1 : boolean;
  signal ptr_deref_2473_store_0_req_0 : boolean;
  signal ptr_deref_2473_store_0_ack_0 : boolean;
  signal ptr_deref_2473_store_0_req_1 : boolean;
  signal ptr_deref_2473_store_0_ack_1 : boolean;
  signal type_cast_2478_inst_req_0 : boolean;
  signal type_cast_2478_inst_ack_0 : boolean;
  signal type_cast_2478_inst_req_1 : boolean;
  signal type_cast_2478_inst_ack_1 : boolean;
  signal if_stmt_2491_branch_req_0 : boolean;
  signal if_stmt_2491_branch_ack_1 : boolean;
  signal if_stmt_2491_branch_ack_0 : boolean;
  signal type_cast_2519_inst_req_0 : boolean;
  signal type_cast_2519_inst_ack_0 : boolean;
  signal type_cast_2519_inst_req_1 : boolean;
  signal type_cast_2519_inst_ack_1 : boolean;
  signal type_cast_2535_inst_req_0 : boolean;
  signal type_cast_2535_inst_ack_0 : boolean;
  signal type_cast_2535_inst_req_1 : boolean;
  signal type_cast_2535_inst_ack_1 : boolean;
  signal if_stmt_2542_branch_req_0 : boolean;
  signal if_stmt_2542_branch_ack_1 : boolean;
  signal if_stmt_2542_branch_ack_0 : boolean;
  signal WPIPE_Block2_done_2578_inst_req_0 : boolean;
  signal WPIPE_Block2_done_2578_inst_ack_0 : boolean;
  signal WPIPE_Block2_done_2578_inst_req_1 : boolean;
  signal WPIPE_Block2_done_2578_inst_ack_1 : boolean;
  signal phi_stmt_2341_req_0 : boolean;
  signal phi_stmt_2348_req_1 : boolean;
  signal phi_stmt_2355_req_1 : boolean;
  signal type_cast_2367_inst_req_0 : boolean;
  signal type_cast_2367_inst_ack_0 : boolean;
  signal type_cast_2367_inst_req_1 : boolean;
  signal type_cast_2367_inst_ack_1 : boolean;
  signal phi_stmt_2362_req_1 : boolean;
  signal type_cast_2347_inst_req_0 : boolean;
  signal type_cast_2347_inst_ack_0 : boolean;
  signal type_cast_2347_inst_req_1 : boolean;
  signal type_cast_2347_inst_ack_1 : boolean;
  signal phi_stmt_2341_req_1 : boolean;
  signal type_cast_2351_inst_req_0 : boolean;
  signal type_cast_2351_inst_ack_0 : boolean;
  signal type_cast_2351_inst_req_1 : boolean;
  signal type_cast_2351_inst_ack_1 : boolean;
  signal phi_stmt_2348_req_0 : boolean;
  signal type_cast_2358_inst_req_0 : boolean;
  signal type_cast_2358_inst_ack_0 : boolean;
  signal type_cast_2358_inst_req_1 : boolean;
  signal type_cast_2358_inst_ack_1 : boolean;
  signal phi_stmt_2355_req_0 : boolean;
  signal type_cast_2365_inst_req_0 : boolean;
  signal type_cast_2365_inst_ack_0 : boolean;
  signal type_cast_2365_inst_req_1 : boolean;
  signal type_cast_2365_inst_ack_1 : boolean;
  signal phi_stmt_2362_req_0 : boolean;
  signal phi_stmt_2341_ack_0 : boolean;
  signal phi_stmt_2348_ack_0 : boolean;
  signal phi_stmt_2355_ack_0 : boolean;
  signal phi_stmt_2362_ack_0 : boolean;
  signal phi_stmt_2549_req_1 : boolean;
  signal type_cast_2559_inst_req_0 : boolean;
  signal type_cast_2559_inst_ack_0 : boolean;
  signal type_cast_2559_inst_req_1 : boolean;
  signal type_cast_2559_inst_ack_1 : boolean;
  signal phi_stmt_2556_req_0 : boolean;
  signal type_cast_2565_inst_req_0 : boolean;
  signal type_cast_2565_inst_ack_0 : boolean;
  signal type_cast_2565_inst_req_1 : boolean;
  signal type_cast_2565_inst_ack_1 : boolean;
  signal phi_stmt_2562_req_0 : boolean;
  signal type_cast_2552_inst_req_0 : boolean;
  signal type_cast_2552_inst_ack_0 : boolean;
  signal type_cast_2552_inst_req_1 : boolean;
  signal type_cast_2552_inst_ack_1 : boolean;
  signal phi_stmt_2549_req_0 : boolean;
  signal type_cast_2561_inst_req_0 : boolean;
  signal type_cast_2561_inst_ack_0 : boolean;
  signal type_cast_2561_inst_req_1 : boolean;
  signal type_cast_2561_inst_ack_1 : boolean;
  signal phi_stmt_2556_req_1 : boolean;
  signal type_cast_2567_inst_req_0 : boolean;
  signal type_cast_2567_inst_ack_0 : boolean;
  signal type_cast_2567_inst_req_1 : boolean;
  signal type_cast_2567_inst_ack_1 : boolean;
  signal phi_stmt_2562_req_1 : boolean;
  signal phi_stmt_2549_ack_0 : boolean;
  signal phi_stmt_2556_ack_0 : boolean;
  signal phi_stmt_2562_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_5768_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5768_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_5768_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5768_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_5768: Block -- control-path 
    signal convTransposeC_CP_5768_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_5768_elements(0) <= convTransposeC_CP_5768_start;
    convTransposeC_CP_5768_symbol <= convTransposeC_CP_5768_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2248_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2248_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2248_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2261_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2261_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2261_update_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2215/$entry
      -- CP-element group 0: 	 branch_block_stmt_2215/branch_block_stmt_2215__entry__
      -- CP-element group 0: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276__entry__
      -- CP-element group 0: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/$entry
      -- CP-element group 0: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2217_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2217_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2217_Sample/rr
      -- 
    cr_5961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(0), ack => type_cast_2248_inst_req_1); -- 
    cr_5989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(0), ack => type_cast_2261_inst_req_1); -- 
    rr_5816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(0), ack => RPIPE_Block2_start_2217_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	92 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2215/merge_stmt_2548__exit__
      -- CP-element group 1: 	 branch_block_stmt_2215/assign_stmt_2574__entry__
      -- CP-element group 1: 	 branch_block_stmt_2215/assign_stmt_2574__exit__
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2215/assign_stmt_2574/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/assign_stmt_2574/$exit
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2362/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2365/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2365/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2365/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2365/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2365/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2365/SplitProtocol/Update/cr
      -- 
    rr_6517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(1), ack => type_cast_2347_inst_req_0); -- 
    cr_6522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(1), ack => type_cast_2347_inst_req_1); -- 
    rr_6540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(1), ack => type_cast_2351_inst_req_0); -- 
    cr_6545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(1), ack => type_cast_2351_inst_req_1); -- 
    rr_6563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(1), ack => type_cast_2358_inst_req_0); -- 
    cr_6568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(1), ack => type_cast_2358_inst_req_1); -- 
    rr_6586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(1), ack => type_cast_2365_inst_req_0); -- 
    cr_6591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(1), ack => type_cast_2365_inst_req_1); -- 
    convTransposeC_CP_5768_elements(1) <= convTransposeC_CP_5768_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2217_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2217_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2217_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2217_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2217_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2217_Update/cr
      -- 
    ra_5817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2217_inst_ack_0, ack => convTransposeC_CP_5768_elements(2)); -- 
    cr_5821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(2), ack => RPIPE_Block2_start_2217_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2217_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2217_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2217_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2220_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2220_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2220_Sample/rr
      -- 
    ca_5822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2217_inst_ack_1, ack => convTransposeC_CP_5768_elements(3)); -- 
    rr_5830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(3), ack => RPIPE_Block2_start_2220_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2220_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2220_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2220_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2220_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2220_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2220_Update/cr
      -- 
    ra_5831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2220_inst_ack_0, ack => convTransposeC_CP_5768_elements(4)); -- 
    cr_5835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(4), ack => RPIPE_Block2_start_2220_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2220_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2220_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2220_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2223_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2223_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2223_Sample/rr
      -- 
    ca_5836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2220_inst_ack_1, ack => convTransposeC_CP_5768_elements(5)); -- 
    rr_5844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(5), ack => RPIPE_Block2_start_2223_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2223_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2223_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2223_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2223_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2223_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2223_Update/$entry
      -- 
    ra_5845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2223_inst_ack_0, ack => convTransposeC_CP_5768_elements(6)); -- 
    cr_5849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(6), ack => RPIPE_Block2_start_2223_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2226_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2226_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2226_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2223_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2223_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2223_update_completed_
      -- 
    ca_5850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2223_inst_ack_1, ack => convTransposeC_CP_5768_elements(7)); -- 
    rr_5858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(7), ack => RPIPE_Block2_start_2226_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2226_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2226_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2226_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2226_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2226_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2226_Update/cr
      -- 
    ra_5859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2226_inst_ack_0, ack => convTransposeC_CP_5768_elements(8)); -- 
    cr_5863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(8), ack => RPIPE_Block2_start_2226_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2226_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2229_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2226_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2226_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2229_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2229_Sample/$entry
      -- 
    ca_5864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2226_inst_ack_1, ack => convTransposeC_CP_5768_elements(9)); -- 
    rr_5872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(9), ack => RPIPE_Block2_start_2229_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2229_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2229_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2229_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2229_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2229_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2229_sample_completed_
      -- 
    ra_5873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2229_inst_ack_0, ack => convTransposeC_CP_5768_elements(10)); -- 
    cr_5877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(10), ack => RPIPE_Block2_start_2229_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2229_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2232_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2232_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2229_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2232_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2229_update_completed_
      -- 
    ca_5878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2229_inst_ack_1, ack => convTransposeC_CP_5768_elements(11)); -- 
    rr_5886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(11), ack => RPIPE_Block2_start_2232_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2232_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2232_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2232_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2232_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2232_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2232_Update/cr
      -- 
    ra_5887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2232_inst_ack_0, ack => convTransposeC_CP_5768_elements(12)); -- 
    cr_5891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(12), ack => RPIPE_Block2_start_2232_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2232_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2235_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2235_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2232_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2232_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2235_sample_start_
      -- 
    ca_5892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2232_inst_ack_1, ack => convTransposeC_CP_5768_elements(13)); -- 
    rr_5900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(13), ack => RPIPE_Block2_start_2235_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2235_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2235_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2235_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2235_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2235_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2235_Update/$entry
      -- 
    ra_5901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2235_inst_ack_0, ack => convTransposeC_CP_5768_elements(14)); -- 
    cr_5905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(14), ack => RPIPE_Block2_start_2235_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2235_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2238_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2235_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2235_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2238_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2238_Sample/$entry
      -- 
    ca_5906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2235_inst_ack_1, ack => convTransposeC_CP_5768_elements(15)); -- 
    rr_5914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(15), ack => RPIPE_Block2_start_2238_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2238_update_start_
      -- CP-element group 16: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2238_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2238_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2238_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2238_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2238_Update/cr
      -- 
    ra_5915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2238_inst_ack_0, ack => convTransposeC_CP_5768_elements(16)); -- 
    cr_5919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(16), ack => RPIPE_Block2_start_2238_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2238_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2241_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2238_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2241_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2238_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2241_sample_start_
      -- 
    ca_5920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2238_inst_ack_1, ack => convTransposeC_CP_5768_elements(17)); -- 
    rr_5928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(17), ack => RPIPE_Block2_start_2241_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2241_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2241_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2241_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2241_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2241_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2241_sample_completed_
      -- 
    ra_5929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2241_inst_ack_0, ack => convTransposeC_CP_5768_elements(18)); -- 
    cr_5933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(18), ack => RPIPE_Block2_start_2241_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2244_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2244_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2241_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2241_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2241_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2244_sample_start_
      -- 
    ca_5934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2241_inst_ack_1, ack => convTransposeC_CP_5768_elements(19)); -- 
    rr_5942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(19), ack => RPIPE_Block2_start_2244_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2244_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2244_update_start_
      -- CP-element group 20: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2244_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2244_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2244_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2244_Update/cr
      -- 
    ra_5943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2244_inst_ack_0, ack => convTransposeC_CP_5768_elements(20)); -- 
    cr_5947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(20), ack => RPIPE_Block2_start_2244_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2257_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2244_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2257_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2257_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2244_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2248_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2244_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2248_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2248_Sample/rr
      -- 
    ca_5948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2244_inst_ack_1, ack => convTransposeC_CP_5768_elements(21)); -- 
    rr_5956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(21), ack => type_cast_2248_inst_req_0); -- 
    rr_5970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(21), ack => RPIPE_Block2_start_2257_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2248_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2248_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2248_Sample/$exit
      -- 
    ra_5957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2248_inst_ack_0, ack => convTransposeC_CP_5768_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2248_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2248_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2248_update_completed_
      -- 
    ca_5962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2248_inst_ack_1, ack => convTransposeC_CP_5768_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2257_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2257_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2257_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2257_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2257_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2257_Update/cr
      -- 
    ra_5971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2257_inst_ack_0, ack => convTransposeC_CP_5768_elements(24)); -- 
    cr_5975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(24), ack => RPIPE_Block2_start_2257_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2269_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2269_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2261_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2257_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2257_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2261_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2257_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2261_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2269_sample_start_
      -- 
    ca_5976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2257_inst_ack_1, ack => convTransposeC_CP_5768_elements(25)); -- 
    rr_5984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(25), ack => type_cast_2261_inst_req_0); -- 
    rr_5998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(25), ack => RPIPE_Block2_start_2269_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2261_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2261_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2261_Sample/ra
      -- 
    ra_5985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2261_inst_ack_0, ack => convTransposeC_CP_5768_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2261_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2261_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/type_cast_2261_Update/$exit
      -- 
    ca_5990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2261_inst_ack_1, ack => convTransposeC_CP_5768_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2269_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2269_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2269_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2269_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2269_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2269_update_start_
      -- 
    ra_5999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2269_inst_ack_0, ack => convTransposeC_CP_5768_elements(28)); -- 
    cr_6003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(28), ack => RPIPE_Block2_start_2269_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2269_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2269_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2269_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2272_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2272_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2272_Sample/$entry
      -- 
    ca_6004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2269_inst_ack_1, ack => convTransposeC_CP_5768_elements(29)); -- 
    rr_6012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(29), ack => RPIPE_Block2_start_2272_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2272_update_start_
      -- CP-element group 30: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2272_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2272_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2272_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2272_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2272_Sample/$exit
      -- 
    ra_6013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2272_inst_ack_0, ack => convTransposeC_CP_5768_elements(30)); -- 
    cr_6017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(30), ack => RPIPE_Block2_start_2272_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2275_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2275_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2275_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2272_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2272_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2272_Update/ca
      -- 
    ca_6018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2272_inst_ack_1, ack => convTransposeC_CP_5768_elements(31)); -- 
    rr_6026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(31), ack => RPIPE_Block2_start_2275_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2275_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2275_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2275_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2275_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2275_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2275_update_start_
      -- 
    ra_6027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2275_inst_ack_0, ack => convTransposeC_CP_5768_elements(32)); -- 
    cr_6031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(32), ack => RPIPE_Block2_start_2275_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2275_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2275_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/RPIPE_Block2_start_2275_update_completed_
      -- 
    ca_6032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2275_inst_ack_1, ack => convTransposeC_CP_5768_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2308_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2312_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2316_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/$entry
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2312_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2312_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2320_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2320_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2316_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2320_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2308_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2320_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2316_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2320_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2320_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2308_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2316_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2312_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2312_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2308_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2316_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2316_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2312_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2308_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2308_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276__exit__
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338__entry__
      -- CP-element group 34: 	 branch_block_stmt_2215/assign_stmt_2218_to_assign_stmt_2276/$exit
      -- 
    cr_6090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(34), ack => type_cast_2320_inst_req_1); -- 
    rr_6085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(34), ack => type_cast_2320_inst_req_0); -- 
    cr_6048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(34), ack => type_cast_2308_inst_req_1); -- 
    cr_6076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(34), ack => type_cast_2316_inst_req_1); -- 
    cr_6062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(34), ack => type_cast_2312_inst_req_1); -- 
    rr_6043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(34), ack => type_cast_2308_inst_req_0); -- 
    rr_6071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(34), ack => type_cast_2316_inst_req_0); -- 
    rr_6057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(34), ack => type_cast_2312_inst_req_0); -- 
    convTransposeC_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(23) & convTransposeC_CP_5768_elements(27) & convTransposeC_CP_5768_elements(33);
      gj_convTransposeC_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2308_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2308_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2308_sample_completed_
      -- 
    ra_6044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2308_inst_ack_0, ack => convTransposeC_CP_5768_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2308_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2308_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2308_update_completed_
      -- 
    ca_6049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2308_inst_ack_1, ack => convTransposeC_CP_5768_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2312_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2312_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2312_Sample/$exit
      -- 
    ra_6058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2312_inst_ack_0, ack => convTransposeC_CP_5768_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2312_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2312_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2312_update_completed_
      -- 
    ca_6063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2312_inst_ack_1, ack => convTransposeC_CP_5768_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2316_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2316_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2316_Sample/ra
      -- 
    ra_6072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2316_inst_ack_0, ack => convTransposeC_CP_5768_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2316_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2316_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2316_Update/ca
      -- 
    ca_6077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2316_inst_ack_1, ack => convTransposeC_CP_5768_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2320_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2320_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2320_sample_completed_
      -- 
    ra_6086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2320_inst_ack_0, ack => convTransposeC_CP_5768_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2320_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2320_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/type_cast_2320_update_completed_
      -- 
    ca_6091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2320_inst_ack_1, ack => convTransposeC_CP_5768_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	82 
    -- CP-element group 43: 	83 
    -- CP-element group 43:  members (18) 
      -- CP-element group 43: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338/$exit
      -- CP-element group 43: 	 branch_block_stmt_2215/assign_stmt_2283_to_assign_stmt_2338__exit__
      -- CP-element group 43: 	 branch_block_stmt_2215/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2341/$entry
      -- CP-element group 43: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2348/$entry
      -- CP-element group 43: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2355/$entry
      -- CP-element group 43: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2362/$entry
      -- CP-element group 43: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2367/$entry
      -- CP-element group 43: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2367/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2367/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2367/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2367/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2367/SplitProtocol/Update/cr
      -- 
    rr_6491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(43), ack => type_cast_2367_inst_req_0); -- 
    cr_6496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(43), ack => type_cast_2367_inst_req_1); -- 
    convTransposeC_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(36) & convTransposeC_CP_5768_elements(38) & convTransposeC_CP_5768_elements(40) & convTransposeC_CP_5768_elements(42);
      gj_convTransposeC_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	104 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2402_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2402_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2402_sample_completed_
      -- 
    ra_6103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2402_inst_ack_0, ack => convTransposeC_CP_5768_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	104 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2402_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2402_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2402_Update/ca
      -- 
    ca_6108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2402_inst_ack_1, ack => convTransposeC_CP_5768_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	104 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2406_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2406_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2406_Sample/ra
      -- 
    ra_6117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2406_inst_ack_0, ack => convTransposeC_CP_5768_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	104 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2406_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2406_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2406_Update/ca
      -- 
    ca_6122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2406_inst_ack_1, ack => convTransposeC_CP_5768_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	104 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2410_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2410_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2410_Sample/ra
      -- 
    ra_6131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2410_inst_ack_0, ack => convTransposeC_CP_5768_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	104 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2410_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2410_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2410_Update/ca
      -- 
    ca_6136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2410_inst_ack_1, ack => convTransposeC_CP_5768_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	104 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2440_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2440_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2440_Sample/ra
      -- 
    ra_6145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2440_inst_ack_0, ack => convTransposeC_CP_5768_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	104 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2440_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2440_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2440_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_final_index_sum_regn_Sample/req
      -- 
    ca_6150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2440_inst_ack_1, ack => convTransposeC_CP_5768_elements(51)); -- 
    req_6175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(51), ack => array_obj_ref_2446_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_final_index_sum_regn_Sample/ack
      -- 
    ack_6176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2446_index_offset_ack_0, ack => convTransposeC_CP_5768_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	104 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2447_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2447_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2447_request/req
      -- 
    ack_6181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2446_index_offset_ack_1, ack => convTransposeC_CP_5768_elements(53)); -- 
    req_6190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(53), ack => addr_of_2447_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2447_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2447_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2447_request/ack
      -- 
    ack_6191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2447_final_reg_ack_0, ack => convTransposeC_CP_5768_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	104 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2447_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2447_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2447_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_Sample/word_access_start/word_0/rr
      -- 
    ack_6196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2447_final_reg_ack_1, ack => convTransposeC_CP_5768_elements(55)); -- 
    rr_6229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(55), ack => ptr_deref_2451_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_Sample/word_access_start/word_0/ra
      -- 
    ra_6230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2451_load_0_ack_0, ack => convTransposeC_CP_5768_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	104 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_Update/ptr_deref_2451_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_Update/ptr_deref_2451_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_Update/ptr_deref_2451_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_Update/ptr_deref_2451_Merge/merge_ack
      -- 
    ca_6241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2451_load_0_ack_1, ack => convTransposeC_CP_5768_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_final_index_sum_regn_Sample/req
      -- 
    req_6271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(58), ack => array_obj_ref_2469_index_offset_req_0); -- 
    convTransposeC_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(45) & convTransposeC_CP_5768_elements(47) & convTransposeC_CP_5768_elements(49);
      gj_convTransposeC_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_final_index_sum_regn_Sample/ack
      -- 
    ack_6272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2469_index_offset_ack_0, ack => convTransposeC_CP_5768_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	104 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2470_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2470_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2470_request/req
      -- 
    ack_6277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2469_index_offset_ack_1, ack => convTransposeC_CP_5768_elements(60)); -- 
    req_6286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(60), ack => addr_of_2470_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2470_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2470_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2470_request/ack
      -- 
    ack_6287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2470_final_reg_ack_0, ack => convTransposeC_CP_5768_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	104 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2470_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2470_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2470_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_word_addrgen/root_register_ack
      -- 
    ack_6292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2470_final_reg_ack_1, ack => convTransposeC_CP_5768_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_Sample/ptr_deref_2473_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_Sample/ptr_deref_2473_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_Sample/ptr_deref_2473_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_Sample/ptr_deref_2473_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_Sample/word_access_start/word_0/rr
      -- 
    rr_6330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(63), ack => ptr_deref_2473_store_0_req_0); -- 
    convTransposeC_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(57) & convTransposeC_CP_5768_elements(62);
      gj_convTransposeC_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_Sample/word_access_start/word_0/ra
      -- 
    ra_6331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2473_store_0_ack_0, ack => convTransposeC_CP_5768_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	104 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_Update/word_access_complete/word_0/ca
      -- 
    ca_6342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2473_store_0_ack_1, ack => convTransposeC_CP_5768_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	104 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2478_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2478_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2478_Sample/ra
      -- 
    ra_6351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2478_inst_ack_0, ack => convTransposeC_CP_5768_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	104 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2478_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2478_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2478_Update/ca
      -- 
    ca_6356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2478_inst_ack_1, ack => convTransposeC_CP_5768_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/$exit
      -- CP-element group 68: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490__exit__
      -- CP-element group 68: 	 branch_block_stmt_2215/if_stmt_2491__entry__
      -- CP-element group 68: 	 branch_block_stmt_2215/if_stmt_2491_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_2215/if_stmt_2491_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_2215/if_stmt_2491_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_2215/if_stmt_2491_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_2215/R_cmp_2492_place
      -- CP-element group 68: 	 branch_block_stmt_2215/if_stmt_2491_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_2215/if_stmt_2491_else_link/$entry
      -- 
    branch_req_6364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(68), ack => if_stmt_2491_branch_req_0); -- 
    convTransposeC_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(52) & convTransposeC_CP_5768_elements(59) & convTransposeC_CP_5768_elements(65) & convTransposeC_CP_5768_elements(67);
      gj_convTransposeC_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	113 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	116 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	119 
    -- CP-element group 69: 	120 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_2215/merge_stmt_2497__exit__
      -- CP-element group 69: 	 branch_block_stmt_2215/assign_stmt_2503__entry__
      -- CP-element group 69: 	 branch_block_stmt_2215/assign_stmt_2503__exit__
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133
      -- CP-element group 69: 	 branch_block_stmt_2215/if_stmt_2491_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_2215/if_stmt_2491_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_2215/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_2215/assign_stmt_2503/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/assign_stmt_2503/$exit
      -- CP-element group 69: 	 branch_block_stmt_2215/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_2215/merge_stmt_2497_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_2215/merge_stmt_2497_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/merge_stmt_2497_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_2215/merge_stmt_2497_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2562/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2567/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2567/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2567/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2567/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2567/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2567/SplitProtocol/Update/cr
      -- 
    if_choice_transition_6369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2491_branch_ack_1, ack => convTransposeC_CP_5768_elements(69)); -- 
    rr_6701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(69), ack => type_cast_2552_inst_req_0); -- 
    cr_6706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(69), ack => type_cast_2552_inst_req_1); -- 
    rr_6724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(69), ack => type_cast_2561_inst_req_0); -- 
    cr_6729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(69), ack => type_cast_2561_inst_req_1); -- 
    rr_6747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(69), ack => type_cast_2567_inst_req_0); -- 
    cr_6752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(69), ack => type_cast_2567_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_2215/merge_stmt_2505__exit__
      -- CP-element group 70: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541__entry__
      -- CP-element group 70: 	 branch_block_stmt_2215/if_stmt_2491_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_2215/if_stmt_2491_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_2215/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/$entry
      -- CP-element group 70: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2519_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2519_update_start_
      -- CP-element group 70: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2519_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2519_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2519_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2519_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2535_update_start_
      -- CP-element group 70: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2535_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2535_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_2215/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_2215/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_2215/merge_stmt_2505_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_2215/merge_stmt_2505_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_2215/merge_stmt_2505_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_2215/merge_stmt_2505_PhiAck/dummy
      -- 
    else_choice_transition_6373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2491_branch_ack_0, ack => convTransposeC_CP_5768_elements(70)); -- 
    rr_6389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(70), ack => type_cast_2519_inst_req_0); -- 
    cr_6394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(70), ack => type_cast_2519_inst_req_1); -- 
    cr_6408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(70), ack => type_cast_2535_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2519_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2519_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2519_Sample/ra
      -- 
    ra_6390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2519_inst_ack_0, ack => convTransposeC_CP_5768_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2519_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2519_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2519_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2535_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2535_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2535_Sample/rr
      -- 
    ca_6395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2519_inst_ack_1, ack => convTransposeC_CP_5768_elements(72)); -- 
    rr_6403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(72), ack => type_cast_2535_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2535_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2535_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2535_Sample/ra
      -- 
    ra_6404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2535_inst_ack_0, ack => convTransposeC_CP_5768_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541__exit__
      -- CP-element group 74: 	 branch_block_stmt_2215/if_stmt_2542__entry__
      -- CP-element group 74: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/$exit
      -- CP-element group 74: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2535_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2535_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2215/assign_stmt_2511_to_assign_stmt_2541/type_cast_2535_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_2215/if_stmt_2542_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2215/if_stmt_2542_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_2215/if_stmt_2542_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_2215/if_stmt_2542_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_2215/R_cmp122_2543_place
      -- CP-element group 74: 	 branch_block_stmt_2215/if_stmt_2542_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2215/if_stmt_2542_else_link/$entry
      -- 
    ca_6409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2535_inst_ack_1, ack => convTransposeC_CP_5768_elements(74)); -- 
    branch_req_6417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(74), ack => if_stmt_2542_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_2215/merge_stmt_2576__exit__
      -- CP-element group 75: 	 branch_block_stmt_2215/assign_stmt_2581__entry__
      -- CP-element group 75: 	 branch_block_stmt_2215/if_stmt_2542_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_2215/if_stmt_2542_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_2215/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_2215/assign_stmt_2581/$entry
      -- CP-element group 75: 	 branch_block_stmt_2215/assign_stmt_2581/WPIPE_Block2_done_2578_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_2215/assign_stmt_2581/WPIPE_Block2_done_2578_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2215/assign_stmt_2581/WPIPE_Block2_done_2578_Sample/req
      -- CP-element group 75: 	 branch_block_stmt_2215/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_2215/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_2215/merge_stmt_2576_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_2215/merge_stmt_2576_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_2215/merge_stmt_2576_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_2215/merge_stmt_2576_PhiAck/dummy
      -- 
    if_choice_transition_6422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2542_branch_ack_1, ack => convTransposeC_CP_5768_elements(75)); -- 
    req_6442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(75), ack => WPIPE_Block2_done_2578_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	105 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	107 
    -- CP-element group 76: 	109 
    -- CP-element group 76: 	110 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_2215/if_stmt_2542_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_2215/if_stmt_2542_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133
      -- CP-element group 76: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/$entry
      -- CP-element group 76: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/$entry
      -- CP-element group 76: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/$entry
      -- CP-element group 76: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2562/$entry
      -- CP-element group 76: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2565/$entry
      -- CP-element group 76: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2565/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2565/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2565/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2565/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2565/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2542_branch_ack_0, ack => convTransposeC_CP_5768_elements(76)); -- 
    rr_6652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(76), ack => type_cast_2559_inst_req_0); -- 
    cr_6657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(76), ack => type_cast_2559_inst_req_1); -- 
    rr_6675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(76), ack => type_cast_2565_inst_req_0); -- 
    cr_6680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(76), ack => type_cast_2565_inst_req_1); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_2215/assign_stmt_2581/WPIPE_Block2_done_2578_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_2215/assign_stmt_2581/WPIPE_Block2_done_2578_update_start_
      -- CP-element group 77: 	 branch_block_stmt_2215/assign_stmt_2581/WPIPE_Block2_done_2578_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_2215/assign_stmt_2581/WPIPE_Block2_done_2578_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_2215/assign_stmt_2581/WPIPE_Block2_done_2578_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_2215/assign_stmt_2581/WPIPE_Block2_done_2578_Update/req
      -- 
    ack_6443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2578_inst_ack_0, ack => convTransposeC_CP_5768_elements(77)); -- 
    req_6447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(77), ack => WPIPE_Block2_done_2578_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_2215/$exit
      -- CP-element group 78: 	 branch_block_stmt_2215/branch_block_stmt_2215__exit__
      -- CP-element group 78: 	 branch_block_stmt_2215/assign_stmt_2581__exit__
      -- CP-element group 78: 	 branch_block_stmt_2215/return__
      -- CP-element group 78: 	 branch_block_stmt_2215/merge_stmt_2583__exit__
      -- CP-element group 78: 	 branch_block_stmt_2215/assign_stmt_2581/$exit
      -- CP-element group 78: 	 branch_block_stmt_2215/assign_stmt_2581/WPIPE_Block2_done_2578_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_2215/assign_stmt_2581/WPIPE_Block2_done_2578_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_2215/assign_stmt_2581/WPIPE_Block2_done_2578_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_2215/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_2215/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_2215/merge_stmt_2583_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_2215/merge_stmt_2583_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_2215/merge_stmt_2583_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_2215/merge_stmt_2583_PhiAck/dummy
      -- 
    ack_6448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2578_inst_ack_1, ack => convTransposeC_CP_5768_elements(78)); -- 
    -- CP-element group 79:  transition  output  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	85 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2341/$exit
      -- CP-element group 79: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2345_konst_delay_trans
      -- CP-element group 79: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_req
      -- 
    phi_stmt_2341_req_6459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2341_req_6459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(79), ack => phi_stmt_2341_req_0); -- 
    -- Element group convTransposeC_CP_5768_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convTransposeC_CP_5768_elements(43), ack => convTransposeC_CP_5768_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  transition  output  delay-element  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	85 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2348/$exit
      -- CP-element group 80: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2354_konst_delay_trans
      -- CP-element group 80: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_req
      -- 
    phi_stmt_2348_req_6467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2348_req_6467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(80), ack => phi_stmt_2348_req_1); -- 
    -- Element group convTransposeC_CP_5768_elements(80) is a control-delay.
    cp_element_80_delay: control_delay_element  generic map(name => " 80_delay", delay_value => 1)  port map(req => convTransposeC_CP_5768_elements(43), ack => convTransposeC_CP_5768_elements(80), clk => clk, reset =>reset);
    -- CP-element group 81:  transition  output  delay-element  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	43 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2355/$exit
      -- CP-element group 81: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2361_konst_delay_trans
      -- CP-element group 81: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_req
      -- 
    phi_stmt_2355_req_6475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2355_req_6475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(81), ack => phi_stmt_2355_req_1); -- 
    -- Element group convTransposeC_CP_5768_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => convTransposeC_CP_5768_elements(43), ack => convTransposeC_CP_5768_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2367/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2367/SplitProtocol/Sample/ra
      -- 
    ra_6492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2367_inst_ack_0, ack => convTransposeC_CP_5768_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	43 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2367/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2367/SplitProtocol/Update/ca
      -- 
    ca_6497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2367_inst_ack_1, ack => convTransposeC_CP_5768_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2362/$exit
      -- CP-element group 84: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2367/$exit
      -- CP-element group 84: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2367/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_req
      -- 
    phi_stmt_2362_req_6498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2362_req_6498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(84), ack => phi_stmt_2362_req_1); -- 
    convTransposeC_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(82) & convTransposeC_CP_5768_elements(83);
      gj_convTransposeC_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	79 
    -- CP-element group 85: 	80 
    -- CP-element group 85: 	81 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	99 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_2215/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(79) & convTransposeC_CP_5768_elements(80) & convTransposeC_CP_5768_elements(81) & convTransposeC_CP_5768_elements(84);
      gj_convTransposeC_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/SplitProtocol/Sample/ra
      -- 
    ra_6518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2347_inst_ack_0, ack => convTransposeC_CP_5768_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/SplitProtocol/Update/ca
      -- 
    ca_6523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2347_inst_ack_1, ack => convTransposeC_CP_5768_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	98 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/$exit
      -- CP-element group 88: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/$exit
      -- CP-element group 88: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/SplitProtocol/$exit
      -- CP-element group 88: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_req
      -- 
    phi_stmt_2341_req_6524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2341_req_6524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(88), ack => phi_stmt_2341_req_1); -- 
    convTransposeC_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(86) & convTransposeC_CP_5768_elements(87);
      gj_convTransposeC_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/SplitProtocol/Sample/ra
      -- 
    ra_6541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2351_inst_ack_0, ack => convTransposeC_CP_5768_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/SplitProtocol/Update/ca
      -- 
    ca_6546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2351_inst_ack_1, ack => convTransposeC_CP_5768_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	98 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/$exit
      -- CP-element group 91: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/$exit
      -- CP-element group 91: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_req
      -- 
    phi_stmt_2348_req_6547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2348_req_6547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(91), ack => phi_stmt_2348_req_0); -- 
    convTransposeC_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(89) & convTransposeC_CP_5768_elements(90);
      gj_convTransposeC_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/SplitProtocol/Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/SplitProtocol/Sample/ra
      -- 
    ra_6564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2358_inst_ack_0, ack => convTransposeC_CP_5768_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/SplitProtocol/Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/SplitProtocol/Update/ca
      -- 
    ca_6569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2358_inst_ack_1, ack => convTransposeC_CP_5768_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	98 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/$exit
      -- CP-element group 94: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/$exit
      -- CP-element group 94: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/SplitProtocol/$exit
      -- CP-element group 94: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_req
      -- 
    phi_stmt_2355_req_6570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2355_req_6570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(94), ack => phi_stmt_2355_req_0); -- 
    convTransposeC_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(92) & convTransposeC_CP_5768_elements(93);
      gj_convTransposeC_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2365/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2365/SplitProtocol/Sample/ra
      -- 
    ra_6587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2365_inst_ack_0, ack => convTransposeC_CP_5768_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2365/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2365/SplitProtocol/Update/ca
      -- 
    ca_6592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2365_inst_ack_1, ack => convTransposeC_CP_5768_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2362/$exit
      -- CP-element group 97: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2365/$exit
      -- CP-element group 97: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_sources/type_cast_2365/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2362/phi_stmt_2362_req
      -- 
    phi_stmt_2362_req_6593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2362_req_6593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(97), ack => phi_stmt_2362_req_0); -- 
    convTransposeC_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(95) & convTransposeC_CP_5768_elements(96);
      gj_convTransposeC_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	88 
    -- CP-element group 98: 	91 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2215/ifx_xend133_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(88) & convTransposeC_CP_5768_elements(91) & convTransposeC_CP_5768_elements(94) & convTransposeC_CP_5768_elements(97);
      gj_convTransposeC_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  merge  fork  transition  place  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	85 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	101 
    -- CP-element group 99: 	102 
    -- CP-element group 99: 	103 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_2215/merge_stmt_2340_PhiReqMerge
      -- CP-element group 99: 	 branch_block_stmt_2215/merge_stmt_2340_PhiAck/$entry
      -- 
    convTransposeC_CP_5768_elements(99) <= OrReduce(convTransposeC_CP_5768_elements(85) & convTransposeC_CP_5768_elements(98));
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_2215/merge_stmt_2340_PhiAck/phi_stmt_2341_ack
      -- 
    phi_stmt_2341_ack_6598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2341_ack_0, ack => convTransposeC_CP_5768_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_2215/merge_stmt_2340_PhiAck/phi_stmt_2348_ack
      -- 
    phi_stmt_2348_ack_6599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2348_ack_0, ack => convTransposeC_CP_5768_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_2215/merge_stmt_2340_PhiAck/phi_stmt_2355_ack
      -- 
    phi_stmt_2355_ack_6600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2355_ack_0, ack => convTransposeC_CP_5768_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	99 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_2215/merge_stmt_2340_PhiAck/phi_stmt_2362_ack
      -- 
    phi_stmt_2362_ack_6601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2362_ack_0, ack => convTransposeC_CP_5768_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  place  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	101 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	44 
    -- CP-element group 104: 	45 
    -- CP-element group 104: 	46 
    -- CP-element group 104: 	47 
    -- CP-element group 104: 	48 
    -- CP-element group 104: 	49 
    -- CP-element group 104: 	50 
    -- CP-element group 104: 	51 
    -- CP-element group 104: 	53 
    -- CP-element group 104: 	55 
    -- CP-element group 104: 	57 
    -- CP-element group 104: 	60 
    -- CP-element group 104: 	62 
    -- CP-element group 104: 	65 
    -- CP-element group 104: 	66 
    -- CP-element group 104: 	67 
    -- CP-element group 104:  members (56) 
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2402_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2402_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/$entry
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2402_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2402_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2402_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2402_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2215/merge_stmt_2340__exit__
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490__entry__
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2406_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2406_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2406_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2406_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2406_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2406_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2410_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2410_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2410_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2410_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2410_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2410_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2440_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2440_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2440_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2440_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2440_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2440_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2447_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2446_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2447_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2447_complete/req
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2451_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2470_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/array_obj_ref_2469_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2470_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/addr_of_2470_complete/req
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/ptr_deref_2473_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2478_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2478_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2478_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2478_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2478_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2215/assign_stmt_2374_to_assign_stmt_2490/type_cast_2478_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2215/merge_stmt_2340_PhiAck/$exit
      -- 
    cr_6107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => type_cast_2402_inst_req_1); -- 
    rr_6102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => type_cast_2402_inst_req_0); -- 
    rr_6116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => type_cast_2406_inst_req_0); -- 
    cr_6121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => type_cast_2406_inst_req_1); -- 
    rr_6130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => type_cast_2410_inst_req_0); -- 
    cr_6135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => type_cast_2410_inst_req_1); -- 
    rr_6144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => type_cast_2440_inst_req_0); -- 
    cr_6149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => type_cast_2440_inst_req_1); -- 
    req_6180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => array_obj_ref_2446_index_offset_req_1); -- 
    req_6195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => addr_of_2447_final_reg_req_1); -- 
    cr_6240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => ptr_deref_2451_load_0_req_1); -- 
    req_6276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => array_obj_ref_2469_index_offset_req_1); -- 
    req_6291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => addr_of_2470_final_reg_req_1); -- 
    cr_6341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => ptr_deref_2473_store_0_req_1); -- 
    rr_6350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => type_cast_2478_inst_req_0); -- 
    cr_6355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => type_cast_2478_inst_req_1); -- 
    convTransposeC_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(100) & convTransposeC_CP_5768_elements(101) & convTransposeC_CP_5768_elements(102) & convTransposeC_CP_5768_elements(103);
      gj_convTransposeC_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  output  delay-element  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	76 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	112 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/$exit
      -- CP-element group 105: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/$exit
      -- CP-element group 105: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2555_konst_delay_trans
      -- CP-element group 105: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_req
      -- 
    phi_stmt_2549_req_6636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2549_req_6636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(105), ack => phi_stmt_2549_req_1); -- 
    -- Element group convTransposeC_CP_5768_elements(105) is a control-delay.
    cp_element_105_delay: control_delay_element  generic map(name => " 105_delay", delay_value => 1)  port map(req => convTransposeC_CP_5768_elements(76), ack => convTransposeC_CP_5768_elements(105), clk => clk, reset =>reset);
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Sample/ra
      -- 
    ra_6653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2559_inst_ack_0, ack => convTransposeC_CP_5768_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	76 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Update/ca
      -- 
    ca_6658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2559_inst_ack_1, ack => convTransposeC_CP_5768_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	112 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/$exit
      -- CP-element group 108: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/$exit
      -- CP-element group 108: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_req
      -- 
    phi_stmt_2556_req_6659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2556_req_6659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(108), ack => phi_stmt_2556_req_0); -- 
    convTransposeC_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(106) & convTransposeC_CP_5768_elements(107);
      gj_convTransposeC_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2565/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2565/SplitProtocol/Sample/ra
      -- 
    ra_6676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2565_inst_ack_0, ack => convTransposeC_CP_5768_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	76 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2565/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2565/SplitProtocol/Update/ca
      -- 
    ca_6681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2565_inst_ack_1, ack => convTransposeC_CP_5768_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2562/$exit
      -- CP-element group 111: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2565/$exit
      -- CP-element group 111: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2565/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_req
      -- 
    phi_stmt_2562_req_6682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2562_req_6682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(111), ack => phi_stmt_2562_req_0); -- 
    convTransposeC_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(109) & convTransposeC_CP_5768_elements(110);
      gj_convTransposeC_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	105 
    -- CP-element group 112: 	108 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	123 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_2215/ifx_xelse_ifx_xend133_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(105) & convTransposeC_CP_5768_elements(108) & convTransposeC_CP_5768_elements(111);
      gj_convTransposeC_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	69 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/SplitProtocol/Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/SplitProtocol/Sample/ra
      -- 
    ra_6702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2552_inst_ack_0, ack => convTransposeC_CP_5768_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/SplitProtocol/Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/SplitProtocol/Update/ca
      -- 
    ca_6707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2552_inst_ack_1, ack => convTransposeC_CP_5768_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	122 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/$exit
      -- CP-element group 115: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/$exit
      -- CP-element group 115: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/SplitProtocol/$exit
      -- CP-element group 115: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_req
      -- 
    phi_stmt_2549_req_6708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2549_req_6708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(115), ack => phi_stmt_2549_req_0); -- 
    convTransposeC_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(113) & convTransposeC_CP_5768_elements(114);
      gj_convTransposeC_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/SplitProtocol/Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/SplitProtocol/Sample/ra
      -- 
    ra_6725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2561_inst_ack_0, ack => convTransposeC_CP_5768_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/SplitProtocol/Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/SplitProtocol/Update/ca
      -- 
    ca_6730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2561_inst_ack_1, ack => convTransposeC_CP_5768_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	122 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/$exit
      -- CP-element group 118: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/$exit
      -- CP-element group 118: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_req
      -- 
    phi_stmt_2556_req_6731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2556_req_6731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(118), ack => phi_stmt_2556_req_1); -- 
    convTransposeC_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(116) & convTransposeC_CP_5768_elements(117);
      gj_convTransposeC_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	69 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2567/SplitProtocol/Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2567/SplitProtocol/Sample/ra
      -- 
    ra_6748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2567_inst_ack_0, ack => convTransposeC_CP_5768_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	69 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2567/SplitProtocol/Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2567/SplitProtocol/Update/ca
      -- 
    ca_6753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2567_inst_ack_1, ack => convTransposeC_CP_5768_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2562/$exit
      -- CP-element group 121: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/$exit
      -- CP-element group 121: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2567/$exit
      -- CP-element group 121: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_sources/type_cast_2567/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2562/phi_stmt_2562_req
      -- 
    phi_stmt_2562_req_6754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2562_req_6754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(121), ack => phi_stmt_2562_req_1); -- 
    convTransposeC_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(119) & convTransposeC_CP_5768_elements(120);
      gj_convTransposeC_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	115 
    -- CP-element group 122: 	118 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2215/ifx_xthen_ifx_xend133_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(115) & convTransposeC_CP_5768_elements(118) & convTransposeC_CP_5768_elements(121);
      gj_convTransposeC_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  fork  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	112 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	126 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_2215/merge_stmt_2548_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_2215/merge_stmt_2548_PhiAck/$entry
      -- 
    convTransposeC_CP_5768_elements(123) <= OrReduce(convTransposeC_CP_5768_elements(112) & convTransposeC_CP_5768_elements(122));
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	127 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_2215/merge_stmt_2548_PhiAck/phi_stmt_2549_ack
      -- 
    phi_stmt_2549_ack_6759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2549_ack_0, ack => convTransposeC_CP_5768_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_2215/merge_stmt_2548_PhiAck/phi_stmt_2556_ack
      -- 
    phi_stmt_2556_ack_6760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2556_ack_0, ack => convTransposeC_CP_5768_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	123 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_2215/merge_stmt_2548_PhiAck/phi_stmt_2562_ack
      -- 
    phi_stmt_2562_ack_6761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2562_ack_0, ack => convTransposeC_CP_5768_elements(126)); -- 
    -- CP-element group 127:  join  transition  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	124 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_2215/merge_stmt_2548_PhiAck/$exit
      -- 
    convTransposeC_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(124) & convTransposeC_CP_5768_elements(125) & convTransposeC_CP_5768_elements(126);
      gj_convTransposeC_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(127), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom86_2468_resized : std_logic_vector(13 downto 0);
    signal R_idxprom86_2468_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2445_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2445_scaled : std_logic_vector(13 downto 0);
    signal add121_2338 : std_logic_vector(31 downto 0);
    signal add45_2289 : std_logic_vector(15 downto 0);
    signal add58_2300 : std_logic_vector(15 downto 0);
    signal add77_2421 : std_logic_vector(63 downto 0);
    signal add79_2431 : std_logic_vector(63 downto 0);
    signal add91_2485 : std_logic_vector(31 downto 0);
    signal add98_2503 : std_logic_vector(15 downto 0);
    signal add_2267 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2379 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2446_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2446_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2446_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2446_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2446_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2446_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2469_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2469_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2469_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2469_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2469_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2469_root_address : std_logic_vector(13 downto 0);
    signal arrayidx82_2448 : std_logic_vector(31 downto 0);
    signal arrayidx87_2471 : std_logic_vector(31 downto 0);
    signal call11_2236 : std_logic_vector(15 downto 0);
    signal call13_2239 : std_logic_vector(15 downto 0);
    signal call14_2242 : std_logic_vector(15 downto 0);
    signal call15_2245 : std_logic_vector(15 downto 0);
    signal call16_2258 : std_logic_vector(15 downto 0);
    signal call18_2270 : std_logic_vector(15 downto 0);
    signal call1_2221 : std_logic_vector(15 downto 0);
    signal call20_2273 : std_logic_vector(15 downto 0);
    signal call22_2276 : std_logic_vector(15 downto 0);
    signal call3_2224 : std_logic_vector(15 downto 0);
    signal call5_2227 : std_logic_vector(15 downto 0);
    signal call7_2230 : std_logic_vector(15 downto 0);
    signal call9_2233 : std_logic_vector(15 downto 0);
    signal call_2218 : std_logic_vector(15 downto 0);
    signal cmp106_2516 : std_logic_vector(0 downto 0);
    signal cmp122_2541 : std_logic_vector(0 downto 0);
    signal cmp_2490 : std_logic_vector(0 downto 0);
    signal conv112_2536 : std_logic_vector(31 downto 0);
    signal conv115_2321 : std_logic_vector(31 downto 0);
    signal conv17_2262 : std_logic_vector(31 downto 0);
    signal conv65_2403 : std_logic_vector(63 downto 0);
    signal conv68_2309 : std_logic_vector(63 downto 0);
    signal conv70_2407 : std_logic_vector(63 downto 0);
    signal conv73_2313 : std_logic_vector(63 downto 0);
    signal conv75_2411 : std_logic_vector(63 downto 0);
    signal conv90_2479 : std_logic_vector(31 downto 0);
    signal conv94_2317 : std_logic_vector(31 downto 0);
    signal conv_2249 : std_logic_vector(31 downto 0);
    signal idxprom86_2464 : std_logic_vector(63 downto 0);
    signal idxprom_2441 : std_logic_vector(63 downto 0);
    signal inc110_2520 : std_logic_vector(15 downto 0);
    signal inc110x_xinput_dim0x_x2_2525 : std_logic_vector(15 downto 0);
    signal inc_2511 : std_logic_vector(15 downto 0);
    signal indvar_2341 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2574 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2562 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_2362 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2556 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2355 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2532 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2549 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2348 : std_logic_vector(15 downto 0);
    signal mul54_2394 : std_logic_vector(15 downto 0);
    signal mul76_2416 : std_logic_vector(63 downto 0);
    signal mul78_2426 : std_logic_vector(63 downto 0);
    signal mul_2384 : std_logic_vector(15 downto 0);
    signal ptr_deref_2451_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2451_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2451_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2451_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2451_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2473_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2473_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2473_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2473_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2473_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2473_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_2255 : std_logic_vector(31 downto 0);
    signal shr116137_2327 : std_logic_vector(31 downto 0);
    signal shr120138_2333 : std_logic_vector(31 downto 0);
    signal shr136_2283 : std_logic_vector(15 downto 0);
    signal shr81_2437 : std_logic_vector(31 downto 0);
    signal shr85_2458 : std_logic_vector(63 downto 0);
    signal sub48_2389 : std_logic_vector(15 downto 0);
    signal sub61_2305 : std_logic_vector(15 downto 0);
    signal sub62_2399 : std_logic_vector(15 downto 0);
    signal sub_2294 : std_logic_vector(15 downto 0);
    signal tmp1_2374 : std_logic_vector(31 downto 0);
    signal tmp83_2452 : std_logic_vector(63 downto 0);
    signal type_cast_2253_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2281_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2287_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2298_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2325_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2331_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2345_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2347_wire : std_logic_vector(31 downto 0);
    signal type_cast_2351_wire : std_logic_vector(15 downto 0);
    signal type_cast_2354_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2358_wire : std_logic_vector(15 downto 0);
    signal type_cast_2361_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2365_wire : std_logic_vector(15 downto 0);
    signal type_cast_2367_wire : std_logic_vector(15 downto 0);
    signal type_cast_2372_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2435_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2456_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2462_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2483_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2501_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2509_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2529_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2552_wire : std_logic_vector(15 downto 0);
    signal type_cast_2555_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2559_wire : std_logic_vector(15 downto 0);
    signal type_cast_2561_wire : std_logic_vector(15 downto 0);
    signal type_cast_2565_wire : std_logic_vector(15 downto 0);
    signal type_cast_2567_wire : std_logic_vector(15 downto 0);
    signal type_cast_2572_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2580_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2446_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2446_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2446_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2446_resized_base_address <= "00000000000000";
    array_obj_ref_2469_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2469_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2469_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2469_resized_base_address <= "00000000000000";
    ptr_deref_2451_word_offset_0 <= "00000000000000";
    ptr_deref_2473_word_offset_0 <= "00000000000000";
    type_cast_2253_wire_constant <= "00000000000000000000000000010000";
    type_cast_2281_wire_constant <= "0000000000000001";
    type_cast_2287_wire_constant <= "1111111111111111";
    type_cast_2298_wire_constant <= "1111111111111111";
    type_cast_2325_wire_constant <= "00000000000000000000000000000010";
    type_cast_2331_wire_constant <= "00000000000000000000000000000001";
    type_cast_2345_wire_constant <= "00000000000000000000000000000000";
    type_cast_2354_wire_constant <= "0000000000000000";
    type_cast_2361_wire_constant <= "0000000000000000";
    type_cast_2372_wire_constant <= "00000000000000000000000000000100";
    type_cast_2435_wire_constant <= "00000000000000000000000000000010";
    type_cast_2456_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2462_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2483_wire_constant <= "00000000000000000000000000000100";
    type_cast_2501_wire_constant <= "0000000000000100";
    type_cast_2509_wire_constant <= "0000000000000001";
    type_cast_2529_wire_constant <= "0000000000000000";
    type_cast_2555_wire_constant <= "0000000000000000";
    type_cast_2572_wire_constant <= "00000000000000000000000000000001";
    type_cast_2580_wire_constant <= "0000000000000001";
    phi_stmt_2341: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2345_wire_constant & type_cast_2347_wire;
      req <= phi_stmt_2341_req_0 & phi_stmt_2341_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2341",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2341_ack_0,
          idata => idata,
          odata => indvar_2341,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2341
    phi_stmt_2348: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2351_wire & type_cast_2354_wire_constant;
      req <= phi_stmt_2348_req_0 & phi_stmt_2348_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2348",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2348_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2348,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2348
    phi_stmt_2355: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2358_wire & type_cast_2361_wire_constant;
      req <= phi_stmt_2355_req_0 & phi_stmt_2355_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2355",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2355_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2355,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2355
    phi_stmt_2362: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2365_wire & type_cast_2367_wire;
      req <= phi_stmt_2362_req_0 & phi_stmt_2362_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2362",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2362_ack_0,
          idata => idata,
          odata => input_dim0x_x2_2362,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2362
    phi_stmt_2549: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2552_wire & type_cast_2555_wire_constant;
      req <= phi_stmt_2549_req_0 & phi_stmt_2549_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2549",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2549_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2549,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2549
    phi_stmt_2556: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2559_wire & type_cast_2561_wire;
      req <= phi_stmt_2556_req_0 & phi_stmt_2556_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2556",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2556_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2556,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2556
    phi_stmt_2562: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2565_wire & type_cast_2567_wire;
      req <= phi_stmt_2562_req_0 & phi_stmt_2562_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2562",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2562_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2562,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2562
    -- flow-through select operator MUX_2531_inst
    input_dim1x_x2_2532 <= type_cast_2529_wire_constant when (cmp106_2516(0) /=  '0') else inc_2511;
    addr_of_2447_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2447_final_reg_req_0;
      addr_of_2447_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2447_final_reg_req_1;
      addr_of_2447_final_reg_ack_1<= rack(0);
      addr_of_2447_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2447_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2446_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_2448,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2470_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2470_final_reg_req_0;
      addr_of_2470_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2470_final_reg_req_1;
      addr_of_2470_final_reg_ack_1<= rack(0);
      addr_of_2470_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2470_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2469_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2471,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2248_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2248_inst_req_0;
      type_cast_2248_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2248_inst_req_1;
      type_cast_2248_inst_ack_1<= rack(0);
      type_cast_2248_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2248_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_2245,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2249,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2261_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2261_inst_req_0;
      type_cast_2261_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2261_inst_req_1;
      type_cast_2261_inst_ack_1<= rack(0);
      type_cast_2261_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2261_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_2258,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_2262,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2308_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2308_inst_req_0;
      type_cast_2308_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2308_inst_req_1;
      type_cast_2308_inst_ack_1<= rack(0);
      type_cast_2308_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2308_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_2276,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_2309,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2312_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2312_inst_req_0;
      type_cast_2312_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2312_inst_req_1;
      type_cast_2312_inst_ack_1<= rack(0);
      type_cast_2312_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2312_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_2273,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2313,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2316_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2316_inst_req_0;
      type_cast_2316_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2316_inst_req_1;
      type_cast_2316_inst_ack_1<= rack(0);
      type_cast_2316_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2316_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2224,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_2317,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2320_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2320_inst_req_0;
      type_cast_2320_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2320_inst_req_1;
      type_cast_2320_inst_ack_1<= rack(0);
      type_cast_2320_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2320_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2218,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_2321,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2347_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2347_inst_req_0;
      type_cast_2347_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2347_inst_req_1;
      type_cast_2347_inst_ack_1<= rack(0);
      type_cast_2347_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2347_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2574,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2347_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2351_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2351_inst_req_0;
      type_cast_2351_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2351_inst_req_1;
      type_cast_2351_inst_ack_1<= rack(0);
      type_cast_2351_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2351_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2549,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2351_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2358_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2358_inst_req_0;
      type_cast_2358_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2358_inst_req_1;
      type_cast_2358_inst_ack_1<= rack(0);
      type_cast_2358_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2358_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2556,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2358_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2365_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2365_inst_req_0;
      type_cast_2365_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2365_inst_req_1;
      type_cast_2365_inst_ack_1<= rack(0);
      type_cast_2365_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2365_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2562,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2365_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2367_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2367_inst_req_0;
      type_cast_2367_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2367_inst_req_1;
      type_cast_2367_inst_ack_1<= rack(0);
      type_cast_2367_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2367_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr136_2283,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2367_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2402_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2402_inst_req_0;
      type_cast_2402_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2402_inst_req_1;
      type_cast_2402_inst_ack_1<= rack(0);
      type_cast_2402_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2402_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2348,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2403,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2406_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2406_inst_req_0;
      type_cast_2406_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2406_inst_req_1;
      type_cast_2406_inst_ack_1<= rack(0);
      type_cast_2406_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2406_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub62_2399,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2407,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2410_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2410_inst_req_0;
      type_cast_2410_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2410_inst_req_1;
      type_cast_2410_inst_ack_1<= rack(0);
      type_cast_2410_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2410_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub48_2389,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2411,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2440_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2440_inst_req_0;
      type_cast_2440_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2440_inst_req_1;
      type_cast_2440_inst_ack_1<= rack(0);
      type_cast_2440_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2440_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr81_2437,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2441,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2478_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2478_inst_req_0;
      type_cast_2478_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2478_inst_req_1;
      type_cast_2478_inst_ack_1<= rack(0);
      type_cast_2478_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2478_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2348,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_2479,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2519_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2519_inst_req_0;
      type_cast_2519_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2519_inst_req_1;
      type_cast_2519_inst_ack_1<= rack(0);
      type_cast_2519_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2519_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp106_2516,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc110_2520,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2535_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2535_inst_req_0;
      type_cast_2535_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2535_inst_req_1;
      type_cast_2535_inst_ack_1<= rack(0);
      type_cast_2535_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2535_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2525,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_2536,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2552_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2552_inst_req_0;
      type_cast_2552_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2552_inst_req_1;
      type_cast_2552_inst_ack_1<= rack(0);
      type_cast_2552_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2552_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add98_2503,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2552_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2559_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2559_inst_req_0;
      type_cast_2559_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2559_inst_req_1;
      type_cast_2559_inst_ack_1<= rack(0);
      type_cast_2559_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2559_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2532,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2559_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2561_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2561_inst_req_0;
      type_cast_2561_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2561_inst_req_1;
      type_cast_2561_inst_ack_1<= rack(0);
      type_cast_2561_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2561_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2355,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2561_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2565_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2565_inst_req_0;
      type_cast_2565_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2565_inst_req_1;
      type_cast_2565_inst_ack_1<= rack(0);
      type_cast_2565_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2565_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2525,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2565_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2567_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2567_inst_req_0;
      type_cast_2567_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2567_inst_req_1;
      type_cast_2567_inst_ack_1<= rack(0);
      type_cast_2567_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2567_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2362,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2567_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2446_index_1_rename
    process(R_idxprom_2445_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2445_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2445_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2446_index_1_resize
    process(idxprom_2441) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2441;
      ov := iv(13 downto 0);
      R_idxprom_2445_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2446_root_address_inst
    process(array_obj_ref_2446_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2446_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2446_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2469_index_1_rename
    process(R_idxprom86_2468_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom86_2468_resized;
      ov(13 downto 0) := iv;
      R_idxprom86_2468_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2469_index_1_resize
    process(idxprom86_2464) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom86_2464;
      ov := iv(13 downto 0);
      R_idxprom86_2468_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2469_root_address_inst
    process(array_obj_ref_2469_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2469_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2469_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2451_addr_0
    process(ptr_deref_2451_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2451_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2451_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2451_base_resize
    process(arrayidx82_2448) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_2448;
      ov := iv(13 downto 0);
      ptr_deref_2451_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2451_gather_scatter
    process(ptr_deref_2451_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2451_data_0;
      ov(63 downto 0) := iv;
      tmp83_2452 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2451_root_address_inst
    process(ptr_deref_2451_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2451_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2451_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2473_addr_0
    process(ptr_deref_2473_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2473_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2473_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2473_base_resize
    process(arrayidx87_2471) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2471;
      ov := iv(13 downto 0);
      ptr_deref_2473_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2473_gather_scatter
    process(tmp83_2452) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp83_2452;
      ov(63 downto 0) := iv;
      ptr_deref_2473_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2473_root_address_inst
    process(ptr_deref_2473_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2473_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2473_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2491_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2490;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2491_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2491_branch_req_0,
          ack0 => if_stmt_2491_branch_ack_0,
          ack1 => if_stmt_2491_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2542_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp122_2541;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2542_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2542_branch_req_0,
          ack0 => if_stmt_2542_branch_ack_0,
          ack1 => if_stmt_2542_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2288_inst
    process(call7_2230) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2230, type_cast_2287_wire_constant, tmp_var);
      add45_2289 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2299_inst
    process(call9_2233) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2233, type_cast_2298_wire_constant, tmp_var);
      add58_2300 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2388_inst
    process(sub_2294, mul_2384) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2294, mul_2384, tmp_var);
      sub48_2389 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2398_inst
    process(sub61_2305, mul54_2394) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub61_2305, mul54_2394, tmp_var);
      sub62_2399 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2502_inst
    process(input_dim2x_x1_2348) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2348, type_cast_2501_wire_constant, tmp_var);
      add98_2503 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2510_inst
    process(input_dim1x_x1_2355) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_2355, type_cast_2509_wire_constant, tmp_var);
      inc_2511 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2524_inst
    process(inc110_2520, input_dim0x_x2_2362) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc110_2520, input_dim0x_x2_2362, tmp_var);
      inc110x_xinput_dim0x_x2_2525 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2337_inst
    process(shr116137_2327, shr120138_2333) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr116137_2327, shr120138_2333, tmp_var);
      add121_2338 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2378_inst
    process(add_2267, tmp1_2374) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_2267, tmp1_2374, tmp_var);
      add_src_0x_x0_2379 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2484_inst
    process(conv90_2479) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv90_2479, type_cast_2483_wire_constant, tmp_var);
      add91_2485 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2573_inst
    process(indvar_2341) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2341, type_cast_2572_wire_constant, tmp_var);
      indvarx_xnext_2574 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2420_inst
    process(mul76_2416, conv70_2407) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul76_2416, conv70_2407, tmp_var);
      add77_2421 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2430_inst
    process(mul78_2426, conv65_2403) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul78_2426, conv65_2403, tmp_var);
      add79_2431 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2463_inst
    process(shr85_2458) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr85_2458, type_cast_2462_wire_constant, tmp_var);
      idxprom86_2464 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2515_inst
    process(inc_2511, call1_2221) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2511, call1_2221, tmp_var);
      cmp106_2516 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2540_inst
    process(conv112_2536, add121_2338) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv112_2536, add121_2338, tmp_var);
      cmp122_2541 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2282_inst
    process(call_2218) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2218, type_cast_2281_wire_constant, tmp_var);
      shr136_2283 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2326_inst
    process(conv115_2321) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_2321, type_cast_2325_wire_constant, tmp_var);
      shr116137_2327 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2332_inst
    process(conv115_2321) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_2321, type_cast_2331_wire_constant, tmp_var);
      shr120138_2333 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2436_inst
    process(add_src_0x_x0_2379) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2379, type_cast_2435_wire_constant, tmp_var);
      shr81_2437 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2457_inst
    process(add79_2431) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_2431, type_cast_2456_wire_constant, tmp_var);
      shr85_2458 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2383_inst
    process(input_dim0x_x2_2362, call13_2239) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_2362, call13_2239, tmp_var);
      mul_2384 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2393_inst
    process(input_dim1x_x1_2355, call13_2239) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2355, call13_2239, tmp_var);
      mul54_2394 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2373_inst
    process(indvar_2341) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2341, type_cast_2372_wire_constant, tmp_var);
      tmp1_2374 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2415_inst
    process(conv75_2411, conv73_2313) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv75_2411, conv73_2313, tmp_var);
      mul76_2416 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2425_inst
    process(add77_2421, conv68_2309) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add77_2421, conv68_2309, tmp_var);
      mul78_2426 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2266_inst
    process(shl_2255, conv17_2262) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2255, conv17_2262, tmp_var);
      add_2267 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2254_inst
    process(conv_2249) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_2249, type_cast_2253_wire_constant, tmp_var);
      shl_2255 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2293_inst
    process(add45_2289, call14_2242) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add45_2289, call14_2242, tmp_var);
      sub_2294 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2304_inst
    process(add58_2300, call14_2242) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add58_2300, call14_2242, tmp_var);
      sub61_2305 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2489_inst
    process(add91_2485, conv94_2317) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add91_2485, conv94_2317, tmp_var);
      cmp_2490 <= tmp_var; --
    end process;
    -- shared split operator group (31) : array_obj_ref_2446_index_offset 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2445_scaled;
      array_obj_ref_2446_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2446_index_offset_req_0;
      array_obj_ref_2446_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2446_index_offset_req_1;
      array_obj_ref_2446_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : array_obj_ref_2469_index_offset 
    ApIntAdd_group_32: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom86_2468_scaled;
      array_obj_ref_2469_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2469_index_offset_req_0;
      array_obj_ref_2469_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2469_index_offset_req_1;
      array_obj_ref_2469_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_32_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared load operator group (0) : ptr_deref_2451_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2451_load_0_req_0;
      ptr_deref_2451_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2451_load_0_req_1;
      ptr_deref_2451_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2451_word_address_0;
      ptr_deref_2451_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2473_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2473_store_0_req_0;
      ptr_deref_2473_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2473_store_0_req_1;
      ptr_deref_2473_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2473_word_address_0;
      data_in <= ptr_deref_2473_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_start_2257_inst RPIPE_Block2_start_2269_inst RPIPE_Block2_start_2272_inst RPIPE_Block2_start_2275_inst RPIPE_Block2_start_2244_inst RPIPE_Block2_start_2241_inst RPIPE_Block2_start_2238_inst RPIPE_Block2_start_2235_inst RPIPE_Block2_start_2232_inst RPIPE_Block2_start_2229_inst RPIPE_Block2_start_2226_inst RPIPE_Block2_start_2223_inst RPIPE_Block2_start_2220_inst RPIPE_Block2_start_2217_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block2_start_2257_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block2_start_2269_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block2_start_2272_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block2_start_2275_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block2_start_2244_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block2_start_2241_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block2_start_2238_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block2_start_2235_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block2_start_2232_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block2_start_2229_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block2_start_2226_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block2_start_2223_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block2_start_2220_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block2_start_2217_inst_req_0;
      RPIPE_Block2_start_2257_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block2_start_2269_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block2_start_2272_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block2_start_2275_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block2_start_2244_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block2_start_2241_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block2_start_2238_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block2_start_2235_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block2_start_2232_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block2_start_2229_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block2_start_2226_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block2_start_2223_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block2_start_2220_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block2_start_2217_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block2_start_2257_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block2_start_2269_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block2_start_2272_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block2_start_2275_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block2_start_2244_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block2_start_2241_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block2_start_2238_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block2_start_2235_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block2_start_2232_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block2_start_2229_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block2_start_2226_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block2_start_2223_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block2_start_2220_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block2_start_2217_inst_req_1;
      RPIPE_Block2_start_2257_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block2_start_2269_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block2_start_2272_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block2_start_2275_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block2_start_2244_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block2_start_2241_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block2_start_2238_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block2_start_2235_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block2_start_2232_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block2_start_2229_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block2_start_2226_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block2_start_2223_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block2_start_2220_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block2_start_2217_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call16_2258 <= data_out(223 downto 208);
      call18_2270 <= data_out(207 downto 192);
      call20_2273 <= data_out(191 downto 176);
      call22_2276 <= data_out(175 downto 160);
      call15_2245 <= data_out(159 downto 144);
      call14_2242 <= data_out(143 downto 128);
      call13_2239 <= data_out(127 downto 112);
      call11_2236 <= data_out(111 downto 96);
      call9_2233 <= data_out(95 downto 80);
      call7_2230 <= data_out(79 downto 64);
      call5_2227 <= data_out(63 downto 48);
      call3_2224 <= data_out(47 downto 32);
      call1_2221 <= data_out(31 downto 16);
      call_2218 <= data_out(15 downto 0);
      Block2_start_read_0_gI: SplitGuardInterface generic map(name => "Block2_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_start_read_0: InputPortRevised -- 
        generic map ( name => "Block2_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_start_pipe_read_req(0),
          oack => Block2_start_pipe_read_ack(0),
          odata => Block2_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2578_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2578_inst_req_0;
      WPIPE_Block2_done_2578_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2578_inst_req_1;
      WPIPE_Block2_done_2578_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2580_wire_constant;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_6778_start: Boolean;
  signal convTransposeD_CP_6778_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block3_start_2647_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2592_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2610_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2592_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2598_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2595_inst_ack_0 : boolean;
  signal type_cast_2620_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2592_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2595_inst_req_0 : boolean;
  signal type_cast_2764_inst_req_1 : boolean;
  signal type_cast_2764_inst_ack_1 : boolean;
  signal type_cast_2699_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2604_inst_req_0 : boolean;
  signal type_cast_2620_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2641_inst_ack_0 : boolean;
  signal type_cast_2691_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2613_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2641_inst_req_0 : boolean;
  signal type_cast_2695_inst_ack_1 : boolean;
  signal type_cast_2772_inst_req_0 : boolean;
  signal type_cast_2772_inst_ack_0 : boolean;
  signal type_cast_2695_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2610_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2601_inst_ack_0 : boolean;
  signal type_cast_2695_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2598_inst_ack_0 : boolean;
  signal type_cast_2633_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2592_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2610_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2641_inst_req_1 : boolean;
  signal type_cast_2699_inst_req_0 : boolean;
  signal type_cast_2691_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2604_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2589_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2610_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2589_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2613_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2647_inst_req_0 : boolean;
  signal type_cast_2764_inst_req_0 : boolean;
  signal type_cast_2764_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2601_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2589_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2641_inst_ack_1 : boolean;
  signal type_cast_2620_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2616_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2629_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2644_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2598_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2595_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2604_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2629_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2601_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2647_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2644_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2613_inst_ack_0 : boolean;
  signal type_cast_2691_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2647_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2613_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2601_inst_ack_1 : boolean;
  signal type_cast_2620_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2644_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2644_inst_ack_0 : boolean;
  signal type_cast_2691_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2589_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2604_inst_ack_1 : boolean;
  signal type_cast_2633_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2595_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2598_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2616_inst_ack_0 : boolean;
  signal type_cast_2772_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2607_inst_ack_1 : boolean;
  signal type_cast_2802_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2607_inst_req_1 : boolean;
  signal type_cast_2802_inst_req_0 : boolean;
  signal type_cast_2802_inst_ack_1 : boolean;
  signal addr_of_2809_final_reg_req_0 : boolean;
  signal addr_of_2809_final_reg_ack_0 : boolean;
  signal addr_of_2809_final_reg_req_1 : boolean;
  signal addr_of_2809_final_reg_ack_1 : boolean;
  signal RPIPE_Block3_start_2607_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2607_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2629_inst_req_1 : boolean;
  signal array_obj_ref_2808_index_offset_ack_0 : boolean;
  signal array_obj_ref_2808_index_offset_req_1 : boolean;
  signal array_obj_ref_2808_index_offset_ack_1 : boolean;
  signal RPIPE_Block3_start_2616_inst_ack_1 : boolean;
  signal type_cast_2695_inst_ack_0 : boolean;
  signal type_cast_2772_inst_ack_1 : boolean;
  signal type_cast_2633_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2616_inst_req_1 : boolean;
  signal type_cast_2633_inst_req_1 : boolean;
  signal type_cast_2768_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2629_inst_ack_1 : boolean;
  signal type_cast_2768_inst_ack_1 : boolean;
  signal type_cast_2699_inst_ack_1 : boolean;
  signal array_obj_ref_2808_index_offset_req_0 : boolean;
  signal type_cast_2768_inst_req_1 : boolean;
  signal type_cast_2699_inst_req_1 : boolean;
  signal type_cast_2768_inst_ack_0 : boolean;
  signal type_cast_2802_inst_ack_0 : boolean;
  signal ptr_deref_2813_load_0_req_0 : boolean;
  signal ptr_deref_2813_load_0_ack_0 : boolean;
  signal ptr_deref_2813_load_0_req_1 : boolean;
  signal ptr_deref_2813_load_0_ack_1 : boolean;
  signal array_obj_ref_2831_index_offset_req_0 : boolean;
  signal array_obj_ref_2831_index_offset_ack_0 : boolean;
  signal array_obj_ref_2831_index_offset_req_1 : boolean;
  signal array_obj_ref_2831_index_offset_ack_1 : boolean;
  signal addr_of_2832_final_reg_req_0 : boolean;
  signal addr_of_2832_final_reg_ack_0 : boolean;
  signal addr_of_2832_final_reg_req_1 : boolean;
  signal addr_of_2832_final_reg_ack_1 : boolean;
  signal ptr_deref_2835_store_0_req_0 : boolean;
  signal ptr_deref_2835_store_0_ack_0 : boolean;
  signal ptr_deref_2835_store_0_req_1 : boolean;
  signal ptr_deref_2835_store_0_ack_1 : boolean;
  signal type_cast_2840_inst_req_0 : boolean;
  signal type_cast_2840_inst_ack_0 : boolean;
  signal type_cast_2840_inst_req_1 : boolean;
  signal type_cast_2840_inst_ack_1 : boolean;
  signal if_stmt_2853_branch_req_0 : boolean;
  signal if_stmt_2853_branch_ack_1 : boolean;
  signal if_stmt_2853_branch_ack_0 : boolean;
  signal type_cast_2881_inst_req_0 : boolean;
  signal type_cast_2881_inst_ack_0 : boolean;
  signal type_cast_2881_inst_req_1 : boolean;
  signal type_cast_2881_inst_ack_1 : boolean;
  signal if_stmt_2900_branch_req_0 : boolean;
  signal if_stmt_2900_branch_ack_1 : boolean;
  signal if_stmt_2900_branch_ack_0 : boolean;
  signal WPIPE_Block3_done_2936_inst_req_0 : boolean;
  signal WPIPE_Block3_done_2936_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_2936_inst_req_1 : boolean;
  signal WPIPE_Block3_done_2936_inst_ack_1 : boolean;
  signal phi_stmt_2703_req_0 : boolean;
  signal phi_stmt_2710_req_0 : boolean;
  signal phi_stmt_2717_req_0 : boolean;
  signal type_cast_2727_inst_req_0 : boolean;
  signal type_cast_2727_inst_ack_0 : boolean;
  signal type_cast_2727_inst_req_1 : boolean;
  signal type_cast_2727_inst_ack_1 : boolean;
  signal phi_stmt_2724_req_0 : boolean;
  signal type_cast_2709_inst_req_0 : boolean;
  signal type_cast_2709_inst_ack_0 : boolean;
  signal type_cast_2709_inst_req_1 : boolean;
  signal type_cast_2709_inst_ack_1 : boolean;
  signal phi_stmt_2703_req_1 : boolean;
  signal type_cast_2716_inst_req_0 : boolean;
  signal type_cast_2716_inst_ack_0 : boolean;
  signal type_cast_2716_inst_req_1 : boolean;
  signal type_cast_2716_inst_ack_1 : boolean;
  signal phi_stmt_2710_req_1 : boolean;
  signal type_cast_2723_inst_req_0 : boolean;
  signal type_cast_2723_inst_ack_0 : boolean;
  signal type_cast_2723_inst_req_1 : boolean;
  signal type_cast_2723_inst_ack_1 : boolean;
  signal phi_stmt_2717_req_1 : boolean;
  signal type_cast_2729_inst_req_0 : boolean;
  signal type_cast_2729_inst_ack_0 : boolean;
  signal type_cast_2729_inst_req_1 : boolean;
  signal type_cast_2729_inst_ack_1 : boolean;
  signal phi_stmt_2724_req_1 : boolean;
  signal phi_stmt_2703_ack_0 : boolean;
  signal phi_stmt_2710_ack_0 : boolean;
  signal phi_stmt_2717_ack_0 : boolean;
  signal phi_stmt_2724_ack_0 : boolean;
  signal phi_stmt_2907_req_1 : boolean;
  signal type_cast_2919_inst_req_0 : boolean;
  signal type_cast_2919_inst_ack_0 : boolean;
  signal type_cast_2919_inst_req_1 : boolean;
  signal type_cast_2919_inst_ack_1 : boolean;
  signal phi_stmt_2914_req_1 : boolean;
  signal type_cast_2925_inst_req_0 : boolean;
  signal type_cast_2925_inst_ack_0 : boolean;
  signal type_cast_2925_inst_req_1 : boolean;
  signal type_cast_2925_inst_ack_1 : boolean;
  signal phi_stmt_2920_req_1 : boolean;
  signal type_cast_2910_inst_req_0 : boolean;
  signal type_cast_2910_inst_ack_0 : boolean;
  signal type_cast_2910_inst_req_1 : boolean;
  signal type_cast_2910_inst_ack_1 : boolean;
  signal phi_stmt_2907_req_0 : boolean;
  signal type_cast_2917_inst_req_0 : boolean;
  signal type_cast_2917_inst_ack_0 : boolean;
  signal type_cast_2917_inst_req_1 : boolean;
  signal type_cast_2917_inst_ack_1 : boolean;
  signal phi_stmt_2914_req_0 : boolean;
  signal type_cast_2923_inst_req_0 : boolean;
  signal type_cast_2923_inst_ack_0 : boolean;
  signal type_cast_2923_inst_req_1 : boolean;
  signal type_cast_2923_inst_ack_1 : boolean;
  signal phi_stmt_2920_req_0 : boolean;
  signal phi_stmt_2907_ack_0 : boolean;
  signal phi_stmt_2914_ack_0 : boolean;
  signal phi_stmt_2920_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_6778_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6778_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_6778_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6778_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_6778: Block -- control-path 
    signal convTransposeD_CP_6778_elements: BooleanArray(123 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_6778_elements(0) <= convTransposeD_CP_6778_start;
    convTransposeD_CP_6778_symbol <= convTransposeD_CP_6778_elements(74);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_2587/branch_block_stmt_2587__entry__
      -- CP-element group 0: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2620_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2620_Update/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2589_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2589_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2633_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2633_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648__entry__
      -- CP-element group 0: 	 branch_block_stmt_2587/$entry
      -- CP-element group 0: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/$entry
      -- CP-element group 0: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2589_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2620_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2633_Update/cr
      -- 
    cr_6971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(0), ack => type_cast_2620_inst_req_1); -- 
    rr_6826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(0), ack => RPIPE_Block3_start_2589_inst_req_0); -- 
    cr_6999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(0), ack => type_cast_2633_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	123 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	82 
    -- CP-element group 1: 	83 
    -- CP-element group 1: 	85 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	88 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	91 
    -- CP-element group 1: 	92 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2587/merge_stmt_2906__exit__
      -- CP-element group 1: 	 branch_block_stmt_2587/assign_stmt_2932__exit__
      -- CP-element group 1: 	 branch_block_stmt_2587/assign_stmt_2932__entry__
      -- CP-element group 1: 	 branch_block_stmt_2587/assign_stmt_2932/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/assign_stmt_2932/$exit
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2723/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2723/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2723/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2723/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2723/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2723/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2724/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2729/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2729/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2729/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2729/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2729/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2729/SplitProtocol/Update/cr
      -- 
    rr_7499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(1), ack => type_cast_2709_inst_req_0); -- 
    cr_7504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(1), ack => type_cast_2709_inst_req_1); -- 
    rr_7522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(1), ack => type_cast_2716_inst_req_0); -- 
    cr_7527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(1), ack => type_cast_2716_inst_req_1); -- 
    rr_7545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(1), ack => type_cast_2723_inst_req_0); -- 
    cr_7550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(1), ack => type_cast_2723_inst_req_1); -- 
    rr_7568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(1), ack => type_cast_2729_inst_req_0); -- 
    cr_7573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(1), ack => type_cast_2729_inst_req_1); -- 
    convTransposeD_CP_6778_elements(1) <= convTransposeD_CP_6778_elements(123);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2589_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2589_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2589_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2589_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2589_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2589_update_start_
      -- 
    ra_6827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2589_inst_ack_0, ack => convTransposeD_CP_6778_elements(2)); -- 
    cr_6831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(2), ack => RPIPE_Block3_start_2589_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2592_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2592_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2592_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2589_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2589_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2589_Update/$exit
      -- 
    ca_6832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2589_inst_ack_1, ack => convTransposeD_CP_6778_elements(3)); -- 
    rr_6840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(3), ack => RPIPE_Block3_start_2592_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2592_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2592_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2592_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2592_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2592_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2592_update_start_
      -- 
    ra_6841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2592_inst_ack_0, ack => convTransposeD_CP_6778_elements(4)); -- 
    cr_6845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(4), ack => RPIPE_Block3_start_2592_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2595_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2595_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2592_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2592_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2592_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2595_Sample/$entry
      -- 
    ca_6846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2592_inst_ack_1, ack => convTransposeD_CP_6778_elements(5)); -- 
    rr_6854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(5), ack => RPIPE_Block3_start_2595_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2595_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2595_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2595_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2595_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2595_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2595_Sample/$exit
      -- 
    ra_6855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2595_inst_ack_0, ack => convTransposeD_CP_6778_elements(6)); -- 
    cr_6859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(6), ack => RPIPE_Block3_start_2595_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2598_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2595_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2595_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2595_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2598_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2598_Sample/rr
      -- 
    ca_6860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2595_inst_ack_1, ack => convTransposeD_CP_6778_elements(7)); -- 
    rr_6868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(7), ack => RPIPE_Block3_start_2598_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2598_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2598_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2598_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2598_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2598_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2598_update_start_
      -- 
    ra_6869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2598_inst_ack_0, ack => convTransposeD_CP_6778_elements(8)); -- 
    cr_6873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(8), ack => RPIPE_Block3_start_2598_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2598_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2598_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2601_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2601_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2598_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2601_sample_start_
      -- 
    ca_6874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2598_inst_ack_1, ack => convTransposeD_CP_6778_elements(9)); -- 
    rr_6882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(9), ack => RPIPE_Block3_start_2601_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2601_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2601_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2601_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2601_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2601_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2601_Update/cr
      -- 
    ra_6883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2601_inst_ack_0, ack => convTransposeD_CP_6778_elements(10)); -- 
    cr_6887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(10), ack => RPIPE_Block3_start_2601_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2601_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2604_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2604_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2601_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2604_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2601_Update/ca
      -- 
    ca_6888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2601_inst_ack_1, ack => convTransposeD_CP_6778_elements(11)); -- 
    rr_6896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(11), ack => RPIPE_Block3_start_2604_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2604_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2604_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2604_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2604_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2604_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2604_Update/cr
      -- 
    ra_6897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2604_inst_ack_0, ack => convTransposeD_CP_6778_elements(12)); -- 
    cr_6901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(12), ack => RPIPE_Block3_start_2604_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2607_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2604_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2604_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2604_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2607_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2607_Sample/$entry
      -- 
    ca_6902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2604_inst_ack_1, ack => convTransposeD_CP_6778_elements(13)); -- 
    rr_6910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(13), ack => RPIPE_Block3_start_2607_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2607_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2607_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2607_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2607_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2607_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2607_sample_completed_
      -- 
    ra_6911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2607_inst_ack_0, ack => convTransposeD_CP_6778_elements(14)); -- 
    cr_6915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(14), ack => RPIPE_Block3_start_2607_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2610_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2610_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2610_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2607_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2607_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2607_update_completed_
      -- 
    ca_6916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2607_inst_ack_1, ack => convTransposeD_CP_6778_elements(15)); -- 
    rr_6924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(15), ack => RPIPE_Block3_start_2610_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2610_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2610_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2610_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2610_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2610_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2610_update_start_
      -- 
    ra_6925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2610_inst_ack_0, ack => convTransposeD_CP_6778_elements(16)); -- 
    cr_6929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(16), ack => RPIPE_Block3_start_2610_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2613_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2610_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2610_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2613_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2610_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2613_Sample/$entry
      -- 
    ca_6930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2610_inst_ack_1, ack => convTransposeD_CP_6778_elements(17)); -- 
    rr_6938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(17), ack => RPIPE_Block3_start_2613_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2613_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2613_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2613_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2613_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2613_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2613_Sample/$exit
      -- 
    ra_6939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2613_inst_ack_0, ack => convTransposeD_CP_6778_elements(18)); -- 
    cr_6943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(18), ack => RPIPE_Block3_start_2613_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2616_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2616_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2616_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2613_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2613_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2613_Update/$exit
      -- 
    ca_6944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2613_inst_ack_1, ack => convTransposeD_CP_6778_elements(19)); -- 
    rr_6952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(19), ack => RPIPE_Block3_start_2616_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2616_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2616_update_start_
      -- CP-element group 20: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2616_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2616_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2616_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2616_Update/cr
      -- 
    ra_6953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2616_inst_ack_0, ack => convTransposeD_CP_6778_elements(20)); -- 
    cr_6957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(20), ack => RPIPE_Block3_start_2616_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2620_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2620_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2616_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2629_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2629_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2629_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2620_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2616_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2616_Update/$exit
      -- 
    ca_6958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2616_inst_ack_1, ack => convTransposeD_CP_6778_elements(21)); -- 
    rr_6966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(21), ack => type_cast_2620_inst_req_0); -- 
    rr_6980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(21), ack => RPIPE_Block3_start_2629_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2620_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2620_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2620_sample_completed_
      -- 
    ra_6967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2620_inst_ack_0, ack => convTransposeD_CP_6778_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2620_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2620_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2620_update_completed_
      -- 
    ca_6972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2620_inst_ack_1, ack => convTransposeD_CP_6778_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2629_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2629_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2629_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2629_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2629_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2629_Update/cr
      -- 
    ra_6981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2629_inst_ack_0, ack => convTransposeD_CP_6778_elements(24)); -- 
    cr_6985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(24), ack => RPIPE_Block3_start_2629_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2629_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2641_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2633_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2633_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2629_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2641_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2641_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2633_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2629_Update/ca
      -- 
    ca_6986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2629_inst_ack_1, ack => convTransposeD_CP_6778_elements(25)); -- 
    rr_6994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(25), ack => type_cast_2633_inst_req_0); -- 
    rr_7008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(25), ack => RPIPE_Block3_start_2641_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2633_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2633_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2633_Sample/$exit
      -- 
    ra_6995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2633_inst_ack_0, ack => convTransposeD_CP_6778_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2633_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2633_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/type_cast_2633_Update/ca
      -- 
    ca_7000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2633_inst_ack_1, ack => convTransposeD_CP_6778_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2641_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2641_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2641_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2641_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2641_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2641_sample_completed_
      -- 
    ra_7009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2641_inst_ack_0, ack => convTransposeD_CP_6778_elements(28)); -- 
    cr_7013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(28), ack => RPIPE_Block3_start_2641_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2641_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2641_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2644_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2644_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2644_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2641_update_completed_
      -- 
    ca_7014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2641_inst_ack_1, ack => convTransposeD_CP_6778_elements(29)); -- 
    rr_7022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(29), ack => RPIPE_Block3_start_2644_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2644_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2644_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2644_update_start_
      -- CP-element group 30: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2644_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2644_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2644_Update/$entry
      -- 
    ra_7023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2644_inst_ack_0, ack => convTransposeD_CP_6778_elements(30)); -- 
    cr_7027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(30), ack => RPIPE_Block3_start_2644_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2647_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2647_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2644_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2644_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2647_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2644_Update/$exit
      -- 
    ca_7028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2644_inst_ack_1, ack => convTransposeD_CP_6778_elements(31)); -- 
    rr_7036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(31), ack => RPIPE_Block3_start_2647_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2647_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2647_update_start_
      -- CP-element group 32: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2647_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2647_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2647_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2647_sample_completed_
      -- 
    ra_7037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2647_inst_ack_0, ack => convTransposeD_CP_6778_elements(32)); -- 
    cr_7041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(32), ack => RPIPE_Block3_start_2647_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2647_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2647_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/RPIPE_Block3_start_2647_Update/$exit
      -- 
    ca_7042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2647_inst_ack_1, ack => convTransposeD_CP_6778_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34:  members (22) 
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2695_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2699_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648__exit__
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2699_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2699_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2695_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2695_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2695_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2699_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/$entry
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700__entry__
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2691_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2691_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2691_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2691_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2691_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2691_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2590_to_assign_stmt_2648/$exit
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2695_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2695_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2699_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2699_Update/$entry
      -- 
    cr_7072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(34), ack => type_cast_2695_inst_req_1); -- 
    rr_7067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(34), ack => type_cast_2695_inst_req_0); -- 
    rr_7081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(34), ack => type_cast_2699_inst_req_0); -- 
    cr_7058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(34), ack => type_cast_2691_inst_req_1); -- 
    rr_7053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(34), ack => type_cast_2691_inst_req_0); -- 
    cr_7086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(34), ack => type_cast_2699_inst_req_1); -- 
    convTransposeD_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(23) & convTransposeD_CP_6778_elements(27) & convTransposeD_CP_6778_elements(33);
      gj_convTransposeD_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2691_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2691_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2691_Sample/$exit
      -- 
    ra_7054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2691_inst_ack_0, ack => convTransposeD_CP_6778_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	41 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2691_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2691_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2691_update_completed_
      -- 
    ca_7059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2691_inst_ack_1, ack => convTransposeD_CP_6778_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2695_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2695_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2695_Sample/ra
      -- 
    ra_7068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2695_inst_ack_0, ack => convTransposeD_CP_6778_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2695_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2695_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2695_update_completed_
      -- 
    ca_7073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2695_inst_ack_1, ack => convTransposeD_CP_6778_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2699_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2699_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2699_sample_completed_
      -- 
    ra_7082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2699_inst_ack_0, ack => convTransposeD_CP_6778_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2699_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2699_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/type_cast_2699_Update/$exit
      -- 
    ca_7087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2699_inst_ack_1, ack => convTransposeD_CP_6778_elements(40)); -- 
    -- CP-element group 41:  join  fork  transition  place  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	36 
    -- CP-element group 41: 	38 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	75 
    -- CP-element group 41: 	76 
    -- CP-element group 41: 	77 
    -- CP-element group 41: 	78 
    -- CP-element group 41: 	79 
    -- CP-element group 41:  members (18) 
      -- CP-element group 41: 	 branch_block_stmt_2587/entry_whilex_xbody
      -- CP-element group 41: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700/$exit
      -- CP-element group 41: 	 branch_block_stmt_2587/assign_stmt_2655_to_assign_stmt_2700__exit__
      -- CP-element group 41: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 41: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2703/$entry
      -- CP-element group 41: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2710/$entry
      -- CP-element group 41: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2717/$entry
      -- CP-element group 41: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2724/$entry
      -- CP-element group 41: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2727/$entry
      -- CP-element group 41: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2727/SplitProtocol/$entry
      -- CP-element group 41: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2727/SplitProtocol/Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2727/SplitProtocol/Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2727/SplitProtocol/Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2727/SplitProtocol/Update/cr
      -- 
    rr_7473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(41), ack => type_cast_2727_inst_req_0); -- 
    cr_7478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(41), ack => type_cast_2727_inst_req_1); -- 
    convTransposeD_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(36) & convTransposeD_CP_6778_elements(38) & convTransposeD_CP_6778_elements(40);
      gj_convTransposeD_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	100 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2764_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2764_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2764_Sample/ra
      -- 
    ra_7099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2764_inst_ack_0, ack => convTransposeD_CP_6778_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	100 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	56 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2764_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2764_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2764_Update/$exit
      -- 
    ca_7104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2764_inst_ack_1, ack => convTransposeD_CP_6778_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	100 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2768_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2768_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2768_Sample/ra
      -- 
    ra_7113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2768_inst_ack_0, ack => convTransposeD_CP_6778_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	100 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	56 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2768_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2768_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2768_Update/$exit
      -- 
    ca_7118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2768_inst_ack_1, ack => convTransposeD_CP_6778_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	100 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2772_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2772_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2772_sample_completed_
      -- 
    ra_7127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2772_inst_ack_0, ack => convTransposeD_CP_6778_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	100 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	56 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2772_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2772_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2772_update_completed_
      -- 
    ca_7132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2772_inst_ack_1, ack => convTransposeD_CP_6778_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	100 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2802_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2802_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2802_Sample/ra
      -- 
    ra_7141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2802_inst_ack_0, ack => convTransposeD_CP_6778_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	100 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (16) 
      -- CP-element group 49: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_index_resize_1/index_resize_req
      -- CP-element group 49: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_index_resize_1/index_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2802_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2802_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_index_resized_1
      -- CP-element group 49: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_index_scaled_1
      -- CP-element group 49: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_index_computed_1
      -- CP-element group 49: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_index_resize_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_index_resize_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_index_scale_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_index_scale_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_index_scale_1/scale_rename_req
      -- CP-element group 49: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_index_scale_1/scale_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_final_index_sum_regn_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_final_index_sum_regn_Sample/req
      -- CP-element group 49: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2802_update_completed_
      -- 
    ca_7146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2802_inst_ack_1, ack => convTransposeD_CP_6778_elements(49)); -- 
    req_7171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(49), ack => array_obj_ref_2808_index_offset_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	66 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_final_index_sum_regn_Sample/ack
      -- CP-element group 50: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_final_index_sum_regn_sample_complete
      -- CP-element group 50: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_final_index_sum_regn_Sample/$exit
      -- 
    ack_7172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2808_index_offset_ack_0, ack => convTransposeD_CP_6778_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	100 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (11) 
      -- CP-element group 51: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_offset_calculated
      -- CP-element group 51: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2809_request/$entry
      -- CP-element group 51: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2809_request/req
      -- CP-element group 51: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_base_plus_offset/$entry
      -- CP-element group 51: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_base_plus_offset/$exit
      -- CP-element group 51: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_base_plus_offset/sum_rename_req
      -- CP-element group 51: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_base_plus_offset/sum_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_final_index_sum_regn_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_final_index_sum_regn_Update/ack
      -- CP-element group 51: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2809_sample_start_
      -- 
    ack_7177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2808_index_offset_ack_1, ack => convTransposeD_CP_6778_elements(51)); -- 
    req_7186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(51), ack => addr_of_2809_final_reg_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2809_request/$exit
      -- CP-element group 52: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2809_request/ack
      -- CP-element group 52: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2809_sample_completed_
      -- 
    ack_7187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2809_final_reg_ack_0, ack => convTransposeD_CP_6778_elements(52)); -- 
    -- CP-element group 53:  join  fork  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	100 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (24) 
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2809_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2809_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2809_complete/ack
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_word_addrgen/$entry
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_word_addrgen/$exit
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_word_addrgen/root_register_req
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_word_addrgen/root_register_ack
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_base_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_word_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_base_address_resized
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_base_addr_resize/$entry
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_base_addr_resize/$exit
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_base_addr_resize/base_resize_req
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_base_addr_resize/base_resize_ack
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_Sample/word_access_start/word_0/rr
      -- 
    ack_7192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2809_final_reg_ack_1, ack => convTransposeD_CP_6778_elements(53)); -- 
    rr_7225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(53), ack => ptr_deref_2813_load_0_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_Sample/word_access_start/word_0/ra
      -- 
    ra_7226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2813_load_0_ack_0, ack => convTransposeD_CP_6778_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	100 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	61 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_Update/word_access_complete/word_0/ca
      -- CP-element group 55: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_Update/ptr_deref_2813_Merge/$entry
      -- CP-element group 55: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_Update/ptr_deref_2813_Merge/$exit
      -- CP-element group 55: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_Update/ptr_deref_2813_Merge/merge_req
      -- CP-element group 55: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_Update/ptr_deref_2813_Merge/merge_ack
      -- 
    ca_7237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2813_load_0_ack_1, ack => convTransposeD_CP_6778_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	43 
    -- CP-element group 56: 	45 
    -- CP-element group 56: 	47 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (13) 
      -- CP-element group 56: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_index_scale_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_index_resized_1
      -- CP-element group 56: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_index_scaled_1
      -- CP-element group 56: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_index_computed_1
      -- CP-element group 56: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_index_resize_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_index_resize_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_index_resize_1/index_resize_req
      -- CP-element group 56: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_index_resize_1/index_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_index_scale_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_index_scale_1/scale_rename_req
      -- CP-element group 56: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_index_scale_1/scale_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_final_index_sum_regn_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_final_index_sum_regn_Sample/req
      -- 
    req_7267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(56), ack => array_obj_ref_2831_index_offset_req_0); -- 
    convTransposeD_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(43) & convTransposeD_CP_6778_elements(45) & convTransposeD_CP_6778_elements(47);
      gj_convTransposeD_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	66 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_final_index_sum_regn_sample_complete
      -- CP-element group 57: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_final_index_sum_regn_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_final_index_sum_regn_Sample/ack
      -- 
    ack_7268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2831_index_offset_ack_0, ack => convTransposeD_CP_6778_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	100 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (11) 
      -- CP-element group 58: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2832_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_offset_calculated
      -- CP-element group 58: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_final_index_sum_regn_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_final_index_sum_regn_Update/ack
      -- CP-element group 58: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_base_plus_offset/$entry
      -- CP-element group 58: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_base_plus_offset/$exit
      -- CP-element group 58: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_base_plus_offset/sum_rename_req
      -- CP-element group 58: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_base_plus_offset/sum_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2832_request/$entry
      -- CP-element group 58: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2832_request/req
      -- 
    ack_7273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2831_index_offset_ack_1, ack => convTransposeD_CP_6778_elements(58)); -- 
    req_7282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(58), ack => addr_of_2832_final_reg_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2832_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2832_request/$exit
      -- CP-element group 59: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2832_request/ack
      -- 
    ack_7283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2832_final_reg_ack_0, ack => convTransposeD_CP_6778_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	100 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (19) 
      -- CP-element group 60: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2832_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2832_complete/$exit
      -- CP-element group 60: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2832_complete/ack
      -- CP-element group 60: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_base_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_word_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_base_address_resized
      -- CP-element group 60: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_base_addr_resize/$entry
      -- CP-element group 60: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_base_addr_resize/$exit
      -- CP-element group 60: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_base_addr_resize/base_resize_req
      -- CP-element group 60: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_base_addr_resize/base_resize_ack
      -- CP-element group 60: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_word_addrgen/$entry
      -- CP-element group 60: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_word_addrgen/$exit
      -- CP-element group 60: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_word_addrgen/root_register_req
      -- CP-element group 60: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_word_addrgen/root_register_ack
      -- 
    ack_7288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2832_final_reg_ack_1, ack => convTransposeD_CP_6778_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	55 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (9) 
      -- CP-element group 61: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_Sample/ptr_deref_2835_Split/$entry
      -- CP-element group 61: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_Sample/ptr_deref_2835_Split/$exit
      -- CP-element group 61: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_Sample/ptr_deref_2835_Split/split_req
      -- CP-element group 61: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_Sample/ptr_deref_2835_Split/split_ack
      -- CP-element group 61: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_Sample/word_access_start/$entry
      -- CP-element group 61: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_Sample/word_access_start/word_0/$entry
      -- CP-element group 61: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_Sample/word_access_start/word_0/rr
      -- 
    rr_7326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(61), ack => ptr_deref_2835_store_0_req_0); -- 
    convTransposeD_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(55) & convTransposeD_CP_6778_elements(60);
      gj_convTransposeD_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (5) 
      -- CP-element group 62: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_Sample/word_access_start/$exit
      -- CP-element group 62: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_Sample/word_access_start/word_0/$exit
      -- CP-element group 62: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_Sample/word_access_start/word_0/ra
      -- 
    ra_7327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2835_store_0_ack_0, ack => convTransposeD_CP_6778_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	100 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	66 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_Update/word_access_complete/$exit
      -- CP-element group 63: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_Update/word_access_complete/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_Update/word_access_complete/word_0/ca
      -- 
    ca_7338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2835_store_0_ack_1, ack => convTransposeD_CP_6778_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	100 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2840_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2840_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2840_Sample/ra
      -- 
    ra_7347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2840_inst_ack_0, ack => convTransposeD_CP_6778_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	100 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2840_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2840_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2840_Update/ca
      -- 
    ca_7352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2840_inst_ack_1, ack => convTransposeD_CP_6778_elements(65)); -- 
    -- CP-element group 66:  branch  join  transition  place  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	50 
    -- CP-element group 66: 	57 
    -- CP-element group 66: 	63 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (10) 
      -- CP-element group 66: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/$exit
      -- CP-element group 66: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852__exit__
      -- CP-element group 66: 	 branch_block_stmt_2587/if_stmt_2853__entry__
      -- CP-element group 66: 	 branch_block_stmt_2587/if_stmt_2853_dead_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2587/if_stmt_2853_eval_test/$entry
      -- CP-element group 66: 	 branch_block_stmt_2587/if_stmt_2853_eval_test/$exit
      -- CP-element group 66: 	 branch_block_stmt_2587/if_stmt_2853_eval_test/branch_req
      -- CP-element group 66: 	 branch_block_stmt_2587/R_cmp_2854_place
      -- CP-element group 66: 	 branch_block_stmt_2587/if_stmt_2853_if_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2587/if_stmt_2853_else_link/$entry
      -- 
    branch_req_7360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(66), ack => if_stmt_2853_branch_req_0); -- 
    convTransposeD_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(50) & convTransposeD_CP_6778_elements(57) & convTransposeD_CP_6778_elements(63) & convTransposeD_CP_6778_elements(65);
      gj_convTransposeD_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	109 
    -- CP-element group 67: 	110 
    -- CP-element group 67: 	112 
    -- CP-element group 67: 	113 
    -- CP-element group 67: 	115 
    -- CP-element group 67: 	116 
    -- CP-element group 67:  members (40) 
      -- CP-element group 67: 	 branch_block_stmt_2587/assign_stmt_2865__exit__
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132
      -- CP-element group 67: 	 branch_block_stmt_2587/assign_stmt_2865__entry__
      -- CP-element group 67: 	 branch_block_stmt_2587/merge_stmt_2859__exit__
      -- CP-element group 67: 	 branch_block_stmt_2587/if_stmt_2853_if_link/$exit
      -- CP-element group 67: 	 branch_block_stmt_2587/if_stmt_2853_if_link/if_choice_transition
      -- CP-element group 67: 	 branch_block_stmt_2587/whilex_xbody_ifx_xthen
      -- CP-element group 67: 	 branch_block_stmt_2587/assign_stmt_2865/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/assign_stmt_2865/$exit
      -- CP-element group 67: 	 branch_block_stmt_2587/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_2587/merge_stmt_2859_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_2587/merge_stmt_2859_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/merge_stmt_2859_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_2587/merge_stmt_2859_PhiAck/dummy
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/SplitProtocol/Update/cr
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Update/cr
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2920/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2923/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2923/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2923/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2923/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2923/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2923/SplitProtocol/Update/cr
      -- 
    if_choice_transition_7365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2853_branch_ack_1, ack => convTransposeD_CP_6778_elements(67)); -- 
    rr_7683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(67), ack => type_cast_2910_inst_req_0); -- 
    cr_7688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(67), ack => type_cast_2910_inst_req_1); -- 
    rr_7706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(67), ack => type_cast_2917_inst_req_0); -- 
    cr_7711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(67), ack => type_cast_2917_inst_req_1); -- 
    rr_7729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(67), ack => type_cast_2923_inst_req_0); -- 
    cr_7734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(67), ack => type_cast_2923_inst_req_1); -- 
    -- CP-element group 68:  fork  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (18) 
      -- CP-element group 68: 	 branch_block_stmt_2587/merge_stmt_2867__exit__
      -- CP-element group 68: 	 branch_block_stmt_2587/assign_stmt_2873_to_assign_stmt_2899__entry__
      -- CP-element group 68: 	 branch_block_stmt_2587/if_stmt_2853_else_link/$exit
      -- CP-element group 68: 	 branch_block_stmt_2587/if_stmt_2853_else_link/else_choice_transition
      -- CP-element group 68: 	 branch_block_stmt_2587/whilex_xbody_ifx_xelse
      -- CP-element group 68: 	 branch_block_stmt_2587/assign_stmt_2873_to_assign_stmt_2899/$entry
      -- CP-element group 68: 	 branch_block_stmt_2587/assign_stmt_2873_to_assign_stmt_2899/type_cast_2881_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_2587/assign_stmt_2873_to_assign_stmt_2899/type_cast_2881_update_start_
      -- CP-element group 68: 	 branch_block_stmt_2587/assign_stmt_2873_to_assign_stmt_2899/type_cast_2881_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2587/assign_stmt_2873_to_assign_stmt_2899/type_cast_2881_Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2587/assign_stmt_2873_to_assign_stmt_2899/type_cast_2881_Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2587/assign_stmt_2873_to_assign_stmt_2899/type_cast_2881_Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2587/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_2587/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 68: 	 branch_block_stmt_2587/merge_stmt_2867_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_2587/merge_stmt_2867_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_2587/merge_stmt_2867_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_2587/merge_stmt_2867_PhiAck/dummy
      -- 
    else_choice_transition_7369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2853_branch_ack_0, ack => convTransposeD_CP_6778_elements(68)); -- 
    rr_7385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(68), ack => type_cast_2881_inst_req_0); -- 
    cr_7390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(68), ack => type_cast_2881_inst_req_1); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2587/assign_stmt_2873_to_assign_stmt_2899/type_cast_2881_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_2587/assign_stmt_2873_to_assign_stmt_2899/type_cast_2881_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_2587/assign_stmt_2873_to_assign_stmt_2899/type_cast_2881_Sample/ra
      -- 
    ra_7386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2881_inst_ack_0, ack => convTransposeD_CP_6778_elements(69)); -- 
    -- CP-element group 70:  branch  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (13) 
      -- CP-element group 70: 	 branch_block_stmt_2587/if_stmt_2900__entry__
      -- CP-element group 70: 	 branch_block_stmt_2587/assign_stmt_2873_to_assign_stmt_2899__exit__
      -- CP-element group 70: 	 branch_block_stmt_2587/assign_stmt_2873_to_assign_stmt_2899/$exit
      -- CP-element group 70: 	 branch_block_stmt_2587/assign_stmt_2873_to_assign_stmt_2899/type_cast_2881_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2587/assign_stmt_2873_to_assign_stmt_2899/type_cast_2881_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2587/assign_stmt_2873_to_assign_stmt_2899/type_cast_2881_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_2587/if_stmt_2900_dead_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2587/if_stmt_2900_eval_test/$entry
      -- CP-element group 70: 	 branch_block_stmt_2587/if_stmt_2900_eval_test/$exit
      -- CP-element group 70: 	 branch_block_stmt_2587/if_stmt_2900_eval_test/branch_req
      -- CP-element group 70: 	 branch_block_stmt_2587/R_cmp121_2901_place
      -- CP-element group 70: 	 branch_block_stmt_2587/if_stmt_2900_if_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2587/if_stmt_2900_else_link/$entry
      -- 
    ca_7391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2881_inst_ack_1, ack => convTransposeD_CP_6778_elements(70)); -- 
    branch_req_7399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(70), ack => if_stmt_2900_branch_req_0); -- 
    -- CP-element group 71:  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (15) 
      -- CP-element group 71: 	 branch_block_stmt_2587/assign_stmt_2939__entry__
      -- CP-element group 71: 	 branch_block_stmt_2587/merge_stmt_2934__exit__
      -- CP-element group 71: 	 branch_block_stmt_2587/if_stmt_2900_if_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_2587/if_stmt_2900_if_link/if_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_2587/ifx_xelse_whilex_xend
      -- CP-element group 71: 	 branch_block_stmt_2587/assign_stmt_2939/$entry
      -- CP-element group 71: 	 branch_block_stmt_2587/assign_stmt_2939/WPIPE_Block3_done_2936_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_2587/assign_stmt_2939/WPIPE_Block3_done_2936_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_2587/assign_stmt_2939/WPIPE_Block3_done_2936_Sample/req
      -- CP-element group 71: 	 branch_block_stmt_2587/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_2587/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 71: 	 branch_block_stmt_2587/merge_stmt_2934_PhiReqMerge
      -- CP-element group 71: 	 branch_block_stmt_2587/merge_stmt_2934_PhiAck/$entry
      -- CP-element group 71: 	 branch_block_stmt_2587/merge_stmt_2934_PhiAck/$exit
      -- CP-element group 71: 	 branch_block_stmt_2587/merge_stmt_2934_PhiAck/dummy
      -- 
    if_choice_transition_7404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2900_branch_ack_1, ack => convTransposeD_CP_6778_elements(71)); -- 
    req_7424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(71), ack => WPIPE_Block3_done_2936_inst_req_0); -- 
    -- CP-element group 72:  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	101 
    -- CP-element group 72: 	102 
    -- CP-element group 72: 	103 
    -- CP-element group 72: 	105 
    -- CP-element group 72: 	106 
    -- CP-element group 72:  members (22) 
      -- CP-element group 72: 	 branch_block_stmt_2587/if_stmt_2900_else_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_2587/if_stmt_2900_else_link/else_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132
      -- CP-element group 72: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/$entry
      -- CP-element group 72: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/$entry
      -- CP-element group 72: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/$entry
      -- CP-element group 72: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Update/cr
      -- CP-element group 72: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2920/$entry
      -- CP-element group 72: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2925/$entry
      -- CP-element group 72: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2925/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2925/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2925/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2925/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2925/SplitProtocol/Update/cr
      -- 
    else_choice_transition_7408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2900_branch_ack_0, ack => convTransposeD_CP_6778_elements(72)); -- 
    rr_7634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(72), ack => type_cast_2919_inst_req_0); -- 
    cr_7639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(72), ack => type_cast_2919_inst_req_1); -- 
    rr_7657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(72), ack => type_cast_2925_inst_req_0); -- 
    cr_7662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(72), ack => type_cast_2925_inst_req_1); -- 
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_2587/assign_stmt_2939/WPIPE_Block3_done_2936_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2587/assign_stmt_2939/WPIPE_Block3_done_2936_update_start_
      -- CP-element group 73: 	 branch_block_stmt_2587/assign_stmt_2939/WPIPE_Block3_done_2936_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2587/assign_stmt_2939/WPIPE_Block3_done_2936_Sample/ack
      -- CP-element group 73: 	 branch_block_stmt_2587/assign_stmt_2939/WPIPE_Block3_done_2936_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_2587/assign_stmt_2939/WPIPE_Block3_done_2936_Update/req
      -- 
    ack_7425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2936_inst_ack_0, ack => convTransposeD_CP_6778_elements(73)); -- 
    req_7429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(73), ack => WPIPE_Block3_done_2936_inst_req_1); -- 
    -- CP-element group 74:  transition  place  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (16) 
      -- CP-element group 74: 	 branch_block_stmt_2587/assign_stmt_2939__exit__
      -- CP-element group 74: 	 branch_block_stmt_2587/branch_block_stmt_2587__exit__
      -- CP-element group 74: 	 $exit
      -- CP-element group 74: 	 branch_block_stmt_2587/return__
      -- CP-element group 74: 	 branch_block_stmt_2587/$exit
      -- CP-element group 74: 	 branch_block_stmt_2587/merge_stmt_2941__exit__
      -- CP-element group 74: 	 branch_block_stmt_2587/assign_stmt_2939/$exit
      -- CP-element group 74: 	 branch_block_stmt_2587/assign_stmt_2939/WPIPE_Block3_done_2936_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2587/assign_stmt_2939/WPIPE_Block3_done_2936_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2587/assign_stmt_2939/WPIPE_Block3_done_2936_Update/ack
      -- CP-element group 74: 	 branch_block_stmt_2587/return___PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_2587/return___PhiReq/$exit
      -- CP-element group 74: 	 branch_block_stmt_2587/merge_stmt_2941_PhiReqMerge
      -- CP-element group 74: 	 branch_block_stmt_2587/merge_stmt_2941_PhiAck/$entry
      -- CP-element group 74: 	 branch_block_stmt_2587/merge_stmt_2941_PhiAck/$exit
      -- CP-element group 74: 	 branch_block_stmt_2587/merge_stmt_2941_PhiAck/dummy
      -- 
    ack_7430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2936_inst_ack_1, ack => convTransposeD_CP_6778_elements(74)); -- 
    -- CP-element group 75:  transition  output  delay-element  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	41 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	81 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2703/$exit
      -- CP-element group 75: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/$exit
      -- CP-element group 75: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2707_konst_delay_trans
      -- CP-element group 75: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_req
      -- 
    phi_stmt_2703_req_7441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2703_req_7441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(75), ack => phi_stmt_2703_req_0); -- 
    -- Element group convTransposeD_CP_6778_elements(75) is a control-delay.
    cp_element_75_delay: control_delay_element  generic map(name => " 75_delay", delay_value => 1)  port map(req => convTransposeD_CP_6778_elements(41), ack => convTransposeD_CP_6778_elements(75), clk => clk, reset =>reset);
    -- CP-element group 76:  transition  output  delay-element  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	41 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	81 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2710/$exit
      -- CP-element group 76: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2714_konst_delay_trans
      -- CP-element group 76: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_req
      -- 
    phi_stmt_2710_req_7449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2710_req_7449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(76), ack => phi_stmt_2710_req_0); -- 
    -- Element group convTransposeD_CP_6778_elements(76) is a control-delay.
    cp_element_76_delay: control_delay_element  generic map(name => " 76_delay", delay_value => 1)  port map(req => convTransposeD_CP_6778_elements(41), ack => convTransposeD_CP_6778_elements(76), clk => clk, reset =>reset);
    -- CP-element group 77:  transition  output  delay-element  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	41 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	81 
    -- CP-element group 77:  members (4) 
      -- CP-element group 77: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2717/$exit
      -- CP-element group 77: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2721_konst_delay_trans
      -- CP-element group 77: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_req
      -- 
    phi_stmt_2717_req_7457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2717_req_7457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(77), ack => phi_stmt_2717_req_0); -- 
    -- Element group convTransposeD_CP_6778_elements(77) is a control-delay.
    cp_element_77_delay: control_delay_element  generic map(name => " 77_delay", delay_value => 1)  port map(req => convTransposeD_CP_6778_elements(41), ack => convTransposeD_CP_6778_elements(77), clk => clk, reset =>reset);
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	41 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2727/SplitProtocol/Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2727/SplitProtocol/Sample/ra
      -- 
    ra_7474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2727_inst_ack_0, ack => convTransposeD_CP_6778_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	41 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2727/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2727/SplitProtocol/Update/ca
      -- 
    ca_7479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2727_inst_ack_1, ack => convTransposeD_CP_6778_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2724/$exit
      -- CP-element group 80: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2727/$exit
      -- CP-element group 80: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2727/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_req
      -- 
    phi_stmt_2724_req_7480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2724_req_7480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(80), ack => phi_stmt_2724_req_0); -- 
    convTransposeD_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(78) & convTransposeD_CP_6778_elements(79);
      gj_convTransposeD_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	75 
    -- CP-element group 81: 	76 
    -- CP-element group 81: 	77 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	95 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2587/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(75) & convTransposeD_CP_6778_elements(76) & convTransposeD_CP_6778_elements(77) & convTransposeD_CP_6778_elements(80);
      gj_convTransposeD_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	1 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/SplitProtocol/Sample/ra
      -- 
    ra_7500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2709_inst_ack_0, ack => convTransposeD_CP_6778_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	1 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/SplitProtocol/Update/ca
      -- 
    ca_7505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2709_inst_ack_1, ack => convTransposeD_CP_6778_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	94 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/$exit
      -- CP-element group 84: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/$exit
      -- CP-element group 84: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_req
      -- 
    phi_stmt_2703_req_7506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2703_req_7506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(84), ack => phi_stmt_2703_req_1); -- 
    convTransposeD_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(82) & convTransposeD_CP_6778_elements(83);
      gj_convTransposeD_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	1 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/SplitProtocol/Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/SplitProtocol/Sample/ra
      -- 
    ra_7523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2716_inst_ack_0, ack => convTransposeD_CP_6778_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/SplitProtocol/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/SplitProtocol/Update/ca
      -- 
    ca_7528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2716_inst_ack_1, ack => convTransposeD_CP_6778_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	94 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/$exit
      -- CP-element group 87: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/$exit
      -- CP-element group 87: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/$exit
      -- CP-element group 87: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/SplitProtocol/$exit
      -- CP-element group 87: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_req
      -- 
    phi_stmt_2710_req_7529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2710_req_7529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(87), ack => phi_stmt_2710_req_1); -- 
    convTransposeD_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(85) & convTransposeD_CP_6778_elements(86);
      gj_convTransposeD_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	1 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2723/SplitProtocol/Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2723/SplitProtocol/Sample/ra
      -- 
    ra_7546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2723_inst_ack_0, ack => convTransposeD_CP_6778_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2723/SplitProtocol/Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2723/SplitProtocol/Update/ca
      -- 
    ca_7551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2723_inst_ack_1, ack => convTransposeD_CP_6778_elements(89)); -- 
    -- CP-element group 90:  join  transition  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	94 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/$exit
      -- CP-element group 90: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/$exit
      -- CP-element group 90: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2723/$exit
      -- CP-element group 90: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2723/SplitProtocol/$exit
      -- CP-element group 90: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_req
      -- 
    phi_stmt_2717_req_7552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2717_req_7552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(90), ack => phi_stmt_2717_req_1); -- 
    convTransposeD_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(88) & convTransposeD_CP_6778_elements(89);
      gj_convTransposeD_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2729/SplitProtocol/Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2729/SplitProtocol/Sample/ra
      -- 
    ra_7569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2729_inst_ack_0, ack => convTransposeD_CP_6778_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2729/SplitProtocol/Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2729/SplitProtocol/Update/ca
      -- 
    ca_7574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2729_inst_ack_1, ack => convTransposeD_CP_6778_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2724/$exit
      -- CP-element group 93: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/$exit
      -- CP-element group 93: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2729/$exit
      -- CP-element group 93: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_sources/type_cast_2729/SplitProtocol/$exit
      -- CP-element group 93: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2724/phi_stmt_2724_req
      -- 
    phi_stmt_2724_req_7575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2724_req_7575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(93), ack => phi_stmt_2724_req_1); -- 
    convTransposeD_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(91) & convTransposeD_CP_6778_elements(92);
      gj_convTransposeD_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	84 
    -- CP-element group 94: 	87 
    -- CP-element group 94: 	90 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_2587/ifx_xend132_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(84) & convTransposeD_CP_6778_elements(87) & convTransposeD_CP_6778_elements(90) & convTransposeD_CP_6778_elements(93);
      gj_convTransposeD_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  merge  fork  transition  place  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	81 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	97 
    -- CP-element group 95: 	98 
    -- CP-element group 95: 	99 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2587/merge_stmt_2702_PhiReqMerge
      -- CP-element group 95: 	 branch_block_stmt_2587/merge_stmt_2702_PhiAck/$entry
      -- 
    convTransposeD_CP_6778_elements(95) <= OrReduce(convTransposeD_CP_6778_elements(81) & convTransposeD_CP_6778_elements(94));
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	100 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_2587/merge_stmt_2702_PhiAck/phi_stmt_2703_ack
      -- 
    phi_stmt_2703_ack_7580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2703_ack_0, ack => convTransposeD_CP_6778_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	100 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_2587/merge_stmt_2702_PhiAck/phi_stmt_2710_ack
      -- 
    phi_stmt_2710_ack_7581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2710_ack_0, ack => convTransposeD_CP_6778_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2587/merge_stmt_2702_PhiAck/phi_stmt_2717_ack
      -- 
    phi_stmt_2717_ack_7582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2717_ack_0, ack => convTransposeD_CP_6778_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	95 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_2587/merge_stmt_2702_PhiAck/phi_stmt_2724_ack
      -- 
    phi_stmt_2724_ack_7583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2724_ack_0, ack => convTransposeD_CP_6778_elements(99)); -- 
    -- CP-element group 100:  join  fork  transition  place  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	96 
    -- CP-element group 100: 	97 
    -- CP-element group 100: 	98 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	42 
    -- CP-element group 100: 	43 
    -- CP-element group 100: 	44 
    -- CP-element group 100: 	45 
    -- CP-element group 100: 	46 
    -- CP-element group 100: 	47 
    -- CP-element group 100: 	48 
    -- CP-element group 100: 	49 
    -- CP-element group 100: 	51 
    -- CP-element group 100: 	53 
    -- CP-element group 100: 	55 
    -- CP-element group 100: 	58 
    -- CP-element group 100: 	60 
    -- CP-element group 100: 	63 
    -- CP-element group 100: 	64 
    -- CP-element group 100: 	65 
    -- CP-element group 100:  members (56) 
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2764_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/$entry
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2768_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2772_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2764_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2764_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2772_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2768_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2764_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2764_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2764_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2587/merge_stmt_2702__exit__
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852__entry__
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2772_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2772_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2772_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2802_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2802_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2802_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2802_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2809_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2809_complete/req
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_final_index_sum_regn_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_final_index_sum_regn_Update/req
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2809_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2768_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2768_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2802_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2808_final_index_sum_regn_update_start
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2768_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2768_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2802_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2772_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_Update/word_access_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_Update/word_access_complete/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2813_Update/word_access_complete/word_0/cr
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2832_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_final_index_sum_regn_update_start
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_final_index_sum_regn_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/array_obj_ref_2831_final_index_sum_regn_Update/req
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2832_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/addr_of_2832_complete/req
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_Update/word_access_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_Update/word_access_complete/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/ptr_deref_2835_Update/word_access_complete/word_0/cr
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2840_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2840_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2840_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2840_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2840_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2587/assign_stmt_2736_to_assign_stmt_2852/type_cast_2840_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2587/merge_stmt_2702_PhiAck/$exit
      -- 
    cr_7103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => type_cast_2764_inst_req_1); -- 
    rr_7126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => type_cast_2772_inst_req_0); -- 
    rr_7098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => type_cast_2764_inst_req_0); -- 
    cr_7131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => type_cast_2772_inst_req_1); -- 
    cr_7145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => type_cast_2802_inst_req_1); -- 
    rr_7140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => type_cast_2802_inst_req_0); -- 
    req_7191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => addr_of_2809_final_reg_req_1); -- 
    req_7176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => array_obj_ref_2808_index_offset_req_1); -- 
    rr_7112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => type_cast_2768_inst_req_0); -- 
    cr_7117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => type_cast_2768_inst_req_1); -- 
    cr_7236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => ptr_deref_2813_load_0_req_1); -- 
    req_7272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => array_obj_ref_2831_index_offset_req_1); -- 
    req_7287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => addr_of_2832_final_reg_req_1); -- 
    cr_7337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => ptr_deref_2835_store_0_req_1); -- 
    rr_7346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => type_cast_2840_inst_req_0); -- 
    cr_7351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => type_cast_2840_inst_req_1); -- 
    convTransposeD_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(96) & convTransposeD_CP_6778_elements(97) & convTransposeD_CP_6778_elements(98) & convTransposeD_CP_6778_elements(99);
      gj_convTransposeD_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  output  delay-element  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	72 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	108 
    -- CP-element group 101:  members (4) 
      -- CP-element group 101: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/$exit
      -- CP-element group 101: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/$exit
      -- CP-element group 101: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2913_konst_delay_trans
      -- CP-element group 101: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_req
      -- 
    phi_stmt_2907_req_7618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2907_req_7618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(101), ack => phi_stmt_2907_req_1); -- 
    -- Element group convTransposeD_CP_6778_elements(101) is a control-delay.
    cp_element_101_delay: control_delay_element  generic map(name => " 101_delay", delay_value => 1)  port map(req => convTransposeD_CP_6778_elements(72), ack => convTransposeD_CP_6778_elements(101), clk => clk, reset =>reset);
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	72 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Sample/ra
      -- 
    ra_7635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2919_inst_ack_0, ack => convTransposeD_CP_6778_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	72 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Update/ca
      -- 
    ca_7640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2919_inst_ack_1, ack => convTransposeD_CP_6778_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	108 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/$exit
      -- CP-element group 104: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/$exit
      -- CP-element group 104: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_req
      -- 
    phi_stmt_2914_req_7641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2914_req_7641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(104), ack => phi_stmt_2914_req_1); -- 
    convTransposeD_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(102) & convTransposeD_CP_6778_elements(103);
      gj_convTransposeD_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	72 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2925/SplitProtocol/Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2925/SplitProtocol/Sample/ra
      -- 
    ra_7658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2925_inst_ack_0, ack => convTransposeD_CP_6778_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	72 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2925/SplitProtocol/Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2925/SplitProtocol/Update/ca
      -- 
    ca_7663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2925_inst_ack_1, ack => convTransposeD_CP_6778_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2920/$exit
      -- CP-element group 107: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2925/$exit
      -- CP-element group 107: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2925/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_req
      -- 
    phi_stmt_2920_req_7664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2920_req_7664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(107), ack => phi_stmt_2920_req_1); -- 
    convTransposeD_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(105) & convTransposeD_CP_6778_elements(106);
      gj_convTransposeD_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	101 
    -- CP-element group 108: 	104 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	119 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_2587/ifx_xelse_ifx_xend132_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(101) & convTransposeD_CP_6778_elements(104) & convTransposeD_CP_6778_elements(107);
      gj_convTransposeD_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	67 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/SplitProtocol/Sample/ra
      -- 
    ra_7684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2910_inst_ack_0, ack => convTransposeD_CP_6778_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	67 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/SplitProtocol/Update/ca
      -- 
    ca_7689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2910_inst_ack_1, ack => convTransposeD_CP_6778_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	118 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/$exit
      -- CP-element group 111: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/$exit
      -- CP-element group 111: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_req
      -- 
    phi_stmt_2907_req_7690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2907_req_7690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(111), ack => phi_stmt_2907_req_0); -- 
    convTransposeD_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(109) & convTransposeD_CP_6778_elements(110);
      gj_convTransposeD_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	67 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Sample/ra
      -- 
    ra_7707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2917_inst_ack_0, ack => convTransposeD_CP_6778_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	67 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Update/ca
      -- 
    ca_7712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2917_inst_ack_1, ack => convTransposeD_CP_6778_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	118 
    -- CP-element group 114:  members (5) 
      -- CP-element group 114: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/$exit
      -- CP-element group 114: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/$exit
      -- CP-element group 114: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/$exit
      -- CP-element group 114: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/$exit
      -- CP-element group 114: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_req
      -- 
    phi_stmt_2914_req_7713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2914_req_7713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(114), ack => phi_stmt_2914_req_0); -- 
    convTransposeD_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(112) & convTransposeD_CP_6778_elements(113);
      gj_convTransposeD_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	67 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2923/SplitProtocol/Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2923/SplitProtocol/Sample/ra
      -- 
    ra_7730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2923_inst_ack_0, ack => convTransposeD_CP_6778_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	67 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2923/SplitProtocol/Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2923/SplitProtocol/Update/ca
      -- 
    ca_7735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2923_inst_ack_1, ack => convTransposeD_CP_6778_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2920/$exit
      -- CP-element group 117: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/$exit
      -- CP-element group 117: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2923/$exit
      -- CP-element group 117: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_sources/type_cast_2923/SplitProtocol/$exit
      -- CP-element group 117: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2920/phi_stmt_2920_req
      -- 
    phi_stmt_2920_req_7736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2920_req_7736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(117), ack => phi_stmt_2920_req_0); -- 
    convTransposeD_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(115) & convTransposeD_CP_6778_elements(116);
      gj_convTransposeD_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	111 
    -- CP-element group 118: 	114 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_2587/ifx_xthen_ifx_xend132_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(111) & convTransposeD_CP_6778_elements(114) & convTransposeD_CP_6778_elements(117);
      gj_convTransposeD_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	108 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119: 	121 
    -- CP-element group 119: 	122 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_2587/merge_stmt_2906_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_2587/merge_stmt_2906_PhiAck/$entry
      -- 
    convTransposeD_CP_6778_elements(119) <= OrReduce(convTransposeD_CP_6778_elements(108) & convTransposeD_CP_6778_elements(118));
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	123 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_2587/merge_stmt_2906_PhiAck/phi_stmt_2907_ack
      -- 
    phi_stmt_2907_ack_7741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2907_ack_0, ack => convTransposeD_CP_6778_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_2587/merge_stmt_2906_PhiAck/phi_stmt_2914_ack
      -- 
    phi_stmt_2914_ack_7742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2914_ack_0, ack => convTransposeD_CP_6778_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	119 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2587/merge_stmt_2906_PhiAck/phi_stmt_2920_ack
      -- 
    phi_stmt_2920_ack_7743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2920_ack_0, ack => convTransposeD_CP_6778_elements(122)); -- 
    -- CP-element group 123:  join  transition  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	120 
    -- CP-element group 123: 	121 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	1 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_2587/merge_stmt_2906_PhiAck/$exit
      -- 
    convTransposeD_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(120) & convTransposeD_CP_6778_elements(121) & convTransposeD_CP_6778_elements(122);
      gj_convTransposeD_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(123), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom91_2830_resized : std_logic_vector(13 downto 0);
    signal R_idxprom91_2830_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2807_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2807_scaled : std_logic_vector(13 downto 0);
    signal add103_2865 : std_logic_vector(15 downto 0);
    signal add32_2666 : std_logic_vector(15 downto 0);
    signal add50_2672 : std_logic_vector(15 downto 0);
    signal add63_2683 : std_logic_vector(15 downto 0);
    signal add82_2783 : std_logic_vector(63 downto 0);
    signal add84_2793 : std_logic_vector(63 downto 0);
    signal add96_2847 : std_logic_vector(31 downto 0);
    signal add_2639 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2741 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2808_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2808_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2808_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2808_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2808_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2808_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2831_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2831_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2831_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2831_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2831_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2831_root_address : std_logic_vector(13 downto 0);
    signal arrayidx87_2810 : std_logic_vector(31 downto 0);
    signal arrayidx92_2833 : std_logic_vector(31 downto 0);
    signal call11_2608 : std_logic_vector(15 downto 0);
    signal call13_2611 : std_logic_vector(15 downto 0);
    signal call14_2614 : std_logic_vector(15 downto 0);
    signal call15_2617 : std_logic_vector(15 downto 0);
    signal call16_2630 : std_logic_vector(15 downto 0);
    signal call18_2642 : std_logic_vector(15 downto 0);
    signal call1_2593 : std_logic_vector(15 downto 0);
    signal call20_2645 : std_logic_vector(15 downto 0);
    signal call22_2648 : std_logic_vector(15 downto 0);
    signal call3_2596 : std_logic_vector(15 downto 0);
    signal call5_2599 : std_logic_vector(15 downto 0);
    signal call7_2602 : std_logic_vector(15 downto 0);
    signal call9_2605 : std_logic_vector(15 downto 0);
    signal call_2590 : std_logic_vector(15 downto 0);
    signal cmp111_2878 : std_logic_vector(0 downto 0);
    signal cmp121_2899 : std_logic_vector(0 downto 0);
    signal cmp_2852 : std_logic_vector(0 downto 0);
    signal conv17_2634 : std_logic_vector(31 downto 0);
    signal conv70_2765 : std_logic_vector(63 downto 0);
    signal conv73_2692 : std_logic_vector(63 downto 0);
    signal conv75_2769 : std_logic_vector(63 downto 0);
    signal conv78_2696 : std_logic_vector(63 downto 0);
    signal conv80_2773 : std_logic_vector(63 downto 0);
    signal conv95_2841 : std_logic_vector(31 downto 0);
    signal conv99_2700 : std_logic_vector(31 downto 0);
    signal conv_2621 : std_logic_vector(31 downto 0);
    signal idxprom91_2826 : std_logic_vector(63 downto 0);
    signal idxprom_2803 : std_logic_vector(63 downto 0);
    signal inc115_2882 : std_logic_vector(15 downto 0);
    signal inc115x_xinput_dim0x_x2_2887 : std_logic_vector(15 downto 0);
    signal inc_2873 : std_logic_vector(15 downto 0);
    signal indvar_2703 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2932 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2920 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_2724 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2914 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2717 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2894 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2907 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2710 : std_logic_vector(15 downto 0);
    signal mul59_2756 : std_logic_vector(15 downto 0);
    signal mul81_2778 : std_logic_vector(63 downto 0);
    signal mul83_2788 : std_logic_vector(63 downto 0);
    signal mul_2746 : std_logic_vector(15 downto 0);
    signal ptr_deref_2813_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2813_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2813_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2813_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2813_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2835_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2835_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2835_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2835_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2835_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2835_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_2627 : std_logic_vector(31 downto 0);
    signal shr135_2655 : std_logic_vector(15 downto 0);
    signal shr31136_2661 : std_logic_vector(15 downto 0);
    signal shr86_2799 : std_logic_vector(31 downto 0);
    signal shr90_2820 : std_logic_vector(63 downto 0);
    signal sub53_2751 : std_logic_vector(15 downto 0);
    signal sub66_2688 : std_logic_vector(15 downto 0);
    signal sub67_2761 : std_logic_vector(15 downto 0);
    signal sub_2677 : std_logic_vector(15 downto 0);
    signal tmp1_2736 : std_logic_vector(31 downto 0);
    signal tmp88_2814 : std_logic_vector(63 downto 0);
    signal type_cast_2625_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2653_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2659_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2670_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2681_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2707_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2709_wire : std_logic_vector(31 downto 0);
    signal type_cast_2714_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2716_wire : std_logic_vector(15 downto 0);
    signal type_cast_2721_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2723_wire : std_logic_vector(15 downto 0);
    signal type_cast_2727_wire : std_logic_vector(15 downto 0);
    signal type_cast_2729_wire : std_logic_vector(15 downto 0);
    signal type_cast_2734_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2797_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2818_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2824_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2845_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2863_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2871_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2891_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2910_wire : std_logic_vector(15 downto 0);
    signal type_cast_2913_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2917_wire : std_logic_vector(15 downto 0);
    signal type_cast_2919_wire : std_logic_vector(15 downto 0);
    signal type_cast_2923_wire : std_logic_vector(15 downto 0);
    signal type_cast_2925_wire : std_logic_vector(15 downto 0);
    signal type_cast_2930_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2938_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2808_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2808_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2808_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2808_resized_base_address <= "00000000000000";
    array_obj_ref_2831_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2831_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2831_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2831_resized_base_address <= "00000000000000";
    ptr_deref_2813_word_offset_0 <= "00000000000000";
    ptr_deref_2835_word_offset_0 <= "00000000000000";
    type_cast_2625_wire_constant <= "00000000000000000000000000010000";
    type_cast_2653_wire_constant <= "0000000000000010";
    type_cast_2659_wire_constant <= "0000000000000001";
    type_cast_2670_wire_constant <= "1111111111111111";
    type_cast_2681_wire_constant <= "1111111111111111";
    type_cast_2707_wire_constant <= "00000000000000000000000000000000";
    type_cast_2714_wire_constant <= "0000000000000000";
    type_cast_2721_wire_constant <= "0000000000000000";
    type_cast_2734_wire_constant <= "00000000000000000000000000000100";
    type_cast_2797_wire_constant <= "00000000000000000000000000000010";
    type_cast_2818_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2824_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2845_wire_constant <= "00000000000000000000000000000100";
    type_cast_2863_wire_constant <= "0000000000000100";
    type_cast_2871_wire_constant <= "0000000000000001";
    type_cast_2891_wire_constant <= "0000000000000000";
    type_cast_2913_wire_constant <= "0000000000000000";
    type_cast_2930_wire_constant <= "00000000000000000000000000000001";
    type_cast_2938_wire_constant <= "0000000000000001";
    phi_stmt_2703: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2707_wire_constant & type_cast_2709_wire;
      req <= phi_stmt_2703_req_0 & phi_stmt_2703_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2703",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2703_ack_0,
          idata => idata,
          odata => indvar_2703,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2703
    phi_stmt_2710: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2714_wire_constant & type_cast_2716_wire;
      req <= phi_stmt_2710_req_0 & phi_stmt_2710_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2710",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2710_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2710,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2710
    phi_stmt_2717: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2721_wire_constant & type_cast_2723_wire;
      req <= phi_stmt_2717_req_0 & phi_stmt_2717_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2717",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2717_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2717,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2717
    phi_stmt_2724: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2727_wire & type_cast_2729_wire;
      req <= phi_stmt_2724_req_0 & phi_stmt_2724_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2724",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2724_ack_0,
          idata => idata,
          odata => input_dim0x_x2_2724,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2724
    phi_stmt_2907: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2910_wire & type_cast_2913_wire_constant;
      req <= phi_stmt_2907_req_0 & phi_stmt_2907_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2907",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2907_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2907,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2907
    phi_stmt_2914: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2917_wire & type_cast_2919_wire;
      req <= phi_stmt_2914_req_0 & phi_stmt_2914_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2914",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2914_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2914,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2914
    phi_stmt_2920: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2923_wire & type_cast_2925_wire;
      req <= phi_stmt_2920_req_0 & phi_stmt_2920_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2920",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2920_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2920,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2920
    -- flow-through select operator MUX_2893_inst
    input_dim1x_x2_2894 <= type_cast_2891_wire_constant when (cmp111_2878(0) /=  '0') else inc_2873;
    addr_of_2809_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2809_final_reg_req_0;
      addr_of_2809_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2809_final_reg_req_1;
      addr_of_2809_final_reg_ack_1<= rack(0);
      addr_of_2809_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2809_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2808_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2810,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2832_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2832_final_reg_req_0;
      addr_of_2832_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2832_final_reg_req_1;
      addr_of_2832_final_reg_ack_1<= rack(0);
      addr_of_2832_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2832_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2831_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx92_2833,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2620_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2620_inst_req_0;
      type_cast_2620_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2620_inst_req_1;
      type_cast_2620_inst_ack_1<= rack(0);
      type_cast_2620_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2620_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_2617,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2621,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2633_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2633_inst_req_0;
      type_cast_2633_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2633_inst_req_1;
      type_cast_2633_inst_ack_1<= rack(0);
      type_cast_2633_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2633_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_2630,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_2634,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2691_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2691_inst_req_0;
      type_cast_2691_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2691_inst_req_1;
      type_cast_2691_inst_ack_1<= rack(0);
      type_cast_2691_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2691_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_2648,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2692,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2695_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2695_inst_req_0;
      type_cast_2695_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2695_inst_req_1;
      type_cast_2695_inst_ack_1<= rack(0);
      type_cast_2695_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2695_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_2645,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv78_2696,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2699_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2699_inst_req_0;
      type_cast_2699_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2699_inst_req_1;
      type_cast_2699_inst_ack_1<= rack(0);
      type_cast_2699_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2699_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2596,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv99_2700,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2709_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2709_inst_req_0;
      type_cast_2709_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2709_inst_req_1;
      type_cast_2709_inst_ack_1<= rack(0);
      type_cast_2709_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2709_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2932,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2709_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2716_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2716_inst_req_0;
      type_cast_2716_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2716_inst_req_1;
      type_cast_2716_inst_ack_1<= rack(0);
      type_cast_2716_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2716_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2907,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2716_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2723_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2723_inst_req_0;
      type_cast_2723_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2723_inst_req_1;
      type_cast_2723_inst_ack_1<= rack(0);
      type_cast_2723_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2723_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2914,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2723_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2727_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2727_inst_req_0;
      type_cast_2727_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2727_inst_req_1;
      type_cast_2727_inst_ack_1<= rack(0);
      type_cast_2727_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2727_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add32_2666,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2727_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2729_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2729_inst_req_0;
      type_cast_2729_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2729_inst_req_1;
      type_cast_2729_inst_ack_1<= rack(0);
      type_cast_2729_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2729_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2920,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2729_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2764_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2764_inst_req_0;
      type_cast_2764_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2764_inst_req_1;
      type_cast_2764_inst_ack_1<= rack(0);
      type_cast_2764_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2764_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2710,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2765,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2768_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2768_inst_req_0;
      type_cast_2768_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2768_inst_req_1;
      type_cast_2768_inst_ack_1<= rack(0);
      type_cast_2768_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2768_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub67_2761,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2769,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2772_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2772_inst_req_0;
      type_cast_2772_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2772_inst_req_1;
      type_cast_2772_inst_ack_1<= rack(0);
      type_cast_2772_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2772_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub53_2751,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv80_2773,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2802_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2802_inst_req_0;
      type_cast_2802_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2802_inst_req_1;
      type_cast_2802_inst_ack_1<= rack(0);
      type_cast_2802_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2802_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr86_2799,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2803,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2840_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2840_inst_req_0;
      type_cast_2840_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2840_inst_req_1;
      type_cast_2840_inst_ack_1<= rack(0);
      type_cast_2840_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2840_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2710,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_2841,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2881_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2881_inst_req_0;
      type_cast_2881_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2881_inst_req_1;
      type_cast_2881_inst_ack_1<= rack(0);
      type_cast_2881_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2881_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp111_2878,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc115_2882,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2910_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2910_inst_req_0;
      type_cast_2910_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2910_inst_req_1;
      type_cast_2910_inst_ack_1<= rack(0);
      type_cast_2910_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2910_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add103_2865,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2910_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2917_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2917_inst_req_0;
      type_cast_2917_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2917_inst_req_1;
      type_cast_2917_inst_ack_1<= rack(0);
      type_cast_2917_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2917_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2717,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2917_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2919_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2919_inst_req_0;
      type_cast_2919_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2919_inst_req_1;
      type_cast_2919_inst_ack_1<= rack(0);
      type_cast_2919_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2919_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2894,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2919_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2923_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2923_inst_req_0;
      type_cast_2923_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2923_inst_req_1;
      type_cast_2923_inst_ack_1<= rack(0);
      type_cast_2923_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2923_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2724,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2923_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2925_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2925_inst_req_0;
      type_cast_2925_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2925_inst_req_1;
      type_cast_2925_inst_ack_1<= rack(0);
      type_cast_2925_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2925_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc115x_xinput_dim0x_x2_2887,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2925_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2808_index_1_rename
    process(R_idxprom_2807_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2807_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2807_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2808_index_1_resize
    process(idxprom_2803) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2803;
      ov := iv(13 downto 0);
      R_idxprom_2807_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2808_root_address_inst
    process(array_obj_ref_2808_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2808_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2808_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2831_index_1_rename
    process(R_idxprom91_2830_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom91_2830_resized;
      ov(13 downto 0) := iv;
      R_idxprom91_2830_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2831_index_1_resize
    process(idxprom91_2826) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom91_2826;
      ov := iv(13 downto 0);
      R_idxprom91_2830_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2831_root_address_inst
    process(array_obj_ref_2831_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2831_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2831_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2813_addr_0
    process(ptr_deref_2813_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2813_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2813_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2813_base_resize
    process(arrayidx87_2810) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2810;
      ov := iv(13 downto 0);
      ptr_deref_2813_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2813_gather_scatter
    process(ptr_deref_2813_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2813_data_0;
      ov(63 downto 0) := iv;
      tmp88_2814 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2813_root_address_inst
    process(ptr_deref_2813_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2813_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2813_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2835_addr_0
    process(ptr_deref_2835_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2835_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2835_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2835_base_resize
    process(arrayidx92_2833) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx92_2833;
      ov := iv(13 downto 0);
      ptr_deref_2835_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2835_gather_scatter
    process(tmp88_2814) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp88_2814;
      ov(63 downto 0) := iv;
      ptr_deref_2835_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2835_root_address_inst
    process(ptr_deref_2835_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2835_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2835_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2853_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2852;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2853_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2853_branch_req_0,
          ack0 => if_stmt_2853_branch_ack_0,
          ack1 => if_stmt_2853_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2900_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp121_2899;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2900_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2900_branch_req_0,
          ack0 => if_stmt_2900_branch_ack_0,
          ack1 => if_stmt_2900_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2665_inst
    process(shr135_2655, shr31136_2661) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr135_2655, shr31136_2661, tmp_var);
      add32_2666 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2671_inst
    process(call7_2602) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2602, type_cast_2670_wire_constant, tmp_var);
      add50_2672 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2682_inst
    process(call9_2605) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2605, type_cast_2681_wire_constant, tmp_var);
      add63_2683 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2750_inst
    process(sub_2677, mul_2746) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2677, mul_2746, tmp_var);
      sub53_2751 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2760_inst
    process(sub66_2688, mul59_2756) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub66_2688, mul59_2756, tmp_var);
      sub67_2761 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2864_inst
    process(input_dim2x_x1_2710) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2710, type_cast_2863_wire_constant, tmp_var);
      add103_2865 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2872_inst
    process(input_dim1x_x1_2717) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_2717, type_cast_2871_wire_constant, tmp_var);
      inc_2873 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2886_inst
    process(inc115_2882, input_dim0x_x2_2724) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc115_2882, input_dim0x_x2_2724, tmp_var);
      inc115x_xinput_dim0x_x2_2887 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2740_inst
    process(add_2639, tmp1_2736) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_2639, tmp1_2736, tmp_var);
      add_src_0x_x0_2741 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2846_inst
    process(conv95_2841) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv95_2841, type_cast_2845_wire_constant, tmp_var);
      add96_2847 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2931_inst
    process(indvar_2703) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2703, type_cast_2930_wire_constant, tmp_var);
      indvarx_xnext_2932 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2782_inst
    process(mul81_2778, conv75_2769) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul81_2778, conv75_2769, tmp_var);
      add82_2783 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2792_inst
    process(mul83_2788, conv70_2765) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul83_2788, conv70_2765, tmp_var);
      add84_2793 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2825_inst
    process(shr90_2820) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr90_2820, type_cast_2824_wire_constant, tmp_var);
      idxprom91_2826 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2877_inst
    process(inc_2873, call1_2593) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2873, call1_2593, tmp_var);
      cmp111_2878 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2898_inst
    process(inc115x_xinput_dim0x_x2_2887, call_2590) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc115x_xinput_dim0x_x2_2887, call_2590, tmp_var);
      cmp121_2899 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2654_inst
    process(call_2590) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2590, type_cast_2653_wire_constant, tmp_var);
      shr135_2655 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2660_inst
    process(call_2590) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2590, type_cast_2659_wire_constant, tmp_var);
      shr31136_2661 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2798_inst
    process(add_src_0x_x0_2741) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2741, type_cast_2797_wire_constant, tmp_var);
      shr86_2799 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2819_inst
    process(add84_2793) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add84_2793, type_cast_2818_wire_constant, tmp_var);
      shr90_2820 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2745_inst
    process(input_dim0x_x2_2724, call13_2611) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_2724, call13_2611, tmp_var);
      mul_2746 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2755_inst
    process(input_dim1x_x1_2717, call13_2611) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2717, call13_2611, tmp_var);
      mul59_2756 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2735_inst
    process(indvar_2703) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2703, type_cast_2734_wire_constant, tmp_var);
      tmp1_2736 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2777_inst
    process(conv80_2773, conv78_2696) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv80_2773, conv78_2696, tmp_var);
      mul81_2778 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2787_inst
    process(add82_2783, conv73_2692) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add82_2783, conv73_2692, tmp_var);
      mul83_2788 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2638_inst
    process(shl_2627, conv17_2634) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2627, conv17_2634, tmp_var);
      add_2639 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2626_inst
    process(conv_2621) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_2621, type_cast_2625_wire_constant, tmp_var);
      shl_2627 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2676_inst
    process(add50_2672, call14_2614) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add50_2672, call14_2614, tmp_var);
      sub_2677 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2687_inst
    process(add63_2683, call14_2614) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add63_2683, call14_2614, tmp_var);
      sub66_2688 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2851_inst
    process(add96_2847, conv99_2700) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add96_2847, conv99_2700, tmp_var);
      cmp_2852 <= tmp_var; --
    end process;
    -- shared split operator group (30) : array_obj_ref_2808_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2807_scaled;
      array_obj_ref_2808_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2808_index_offset_req_0;
      array_obj_ref_2808_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2808_index_offset_req_1;
      array_obj_ref_2808_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : array_obj_ref_2831_index_offset 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom91_2830_scaled;
      array_obj_ref_2831_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2831_index_offset_req_0;
      array_obj_ref_2831_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2831_index_offset_req_1;
      array_obj_ref_2831_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared load operator group (0) : ptr_deref_2813_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2813_load_0_req_0;
      ptr_deref_2813_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2813_load_0_req_1;
      ptr_deref_2813_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2813_word_address_0;
      ptr_deref_2813_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2835_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2835_store_0_req_0;
      ptr_deref_2835_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2835_store_0_req_1;
      ptr_deref_2835_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2835_word_address_0;
      data_in <= ptr_deref_2835_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_start_2589_inst RPIPE_Block3_start_2592_inst RPIPE_Block3_start_2595_inst RPIPE_Block3_start_2598_inst RPIPE_Block3_start_2601_inst RPIPE_Block3_start_2604_inst RPIPE_Block3_start_2607_inst RPIPE_Block3_start_2610_inst RPIPE_Block3_start_2613_inst RPIPE_Block3_start_2616_inst RPIPE_Block3_start_2629_inst RPIPE_Block3_start_2641_inst RPIPE_Block3_start_2644_inst RPIPE_Block3_start_2647_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block3_start_2589_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block3_start_2592_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block3_start_2595_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block3_start_2598_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block3_start_2601_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block3_start_2604_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block3_start_2607_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block3_start_2610_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block3_start_2613_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block3_start_2616_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block3_start_2629_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block3_start_2641_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block3_start_2644_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block3_start_2647_inst_req_0;
      RPIPE_Block3_start_2589_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block3_start_2592_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block3_start_2595_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block3_start_2598_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block3_start_2601_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block3_start_2604_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block3_start_2607_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block3_start_2610_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block3_start_2613_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block3_start_2616_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block3_start_2629_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block3_start_2641_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block3_start_2644_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block3_start_2647_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block3_start_2589_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block3_start_2592_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block3_start_2595_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block3_start_2598_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block3_start_2601_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block3_start_2604_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block3_start_2607_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block3_start_2610_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block3_start_2613_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block3_start_2616_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block3_start_2629_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block3_start_2641_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block3_start_2644_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block3_start_2647_inst_req_1;
      RPIPE_Block3_start_2589_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block3_start_2592_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block3_start_2595_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block3_start_2598_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block3_start_2601_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block3_start_2604_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block3_start_2607_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block3_start_2610_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block3_start_2613_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block3_start_2616_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block3_start_2629_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block3_start_2641_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block3_start_2644_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block3_start_2647_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call_2590 <= data_out(223 downto 208);
      call1_2593 <= data_out(207 downto 192);
      call3_2596 <= data_out(191 downto 176);
      call5_2599 <= data_out(175 downto 160);
      call7_2602 <= data_out(159 downto 144);
      call9_2605 <= data_out(143 downto 128);
      call11_2608 <= data_out(127 downto 112);
      call13_2611 <= data_out(111 downto 96);
      call14_2614 <= data_out(95 downto 80);
      call15_2617 <= data_out(79 downto 64);
      call16_2630 <= data_out(63 downto 48);
      call18_2642 <= data_out(47 downto 32);
      call20_2645 <= data_out(31 downto 16);
      call22_2648 <= data_out(15 downto 0);
      Block3_start_read_0_gI: SplitGuardInterface generic map(name => "Block3_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_start_read_0: InputPortRevised -- 
        generic map ( name => "Block3_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_start_pipe_read_req(0),
          oack => Block3_start_pipe_read_ack(0),
          odata => Block3_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_2936_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_2936_inst_req_0;
      WPIPE_Block3_done_2936_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_2936_inst_req_1;
      WPIPE_Block3_done_2936_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2938_wire_constant;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    T : out  std_logic_vector(63 downto 0);
    timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
    timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal T_buffer :  std_logic_vector(63 downto 0);
  signal T_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_timer_resp_34_inst_req_0 : boolean;
  signal RPIPE_timer_resp_34_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_34_inst_req_1 : boolean;
  signal RPIPE_timer_resp_34_inst_ack_1 : boolean;
  signal WPIPE_timer_req_29_inst_req_0 : boolean;
  signal WPIPE_timer_req_29_inst_ack_0 : boolean;
  signal WPIPE_timer_req_29_inst_req_1 : boolean;
  signal WPIPE_timer_req_29_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= T_buffer;
  T <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_sample_start_
      -- CP-element group 0: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Sample/rr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_32_to_assign_stmt_35/$entry
      -- CP-element group 0: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_sample_start_
      -- CP-element group 0: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Sample/req
      -- 
    rr_27_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_27_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => RPIPE_timer_resp_34_inst_req_0); -- 
    req_13_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_13_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => WPIPE_timer_req_29_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_sample_completed_
      -- CP-element group 1: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_update_start_
      -- CP-element group 1: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Sample/ack
      -- CP-element group 1: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Update/$entry
      -- CP-element group 1: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Update/req
      -- 
    ack_14_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_29_inst_ack_0, ack => timer_CP_0_elements(1)); -- 
    req_18_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_18_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(1), ack => WPIPE_timer_req_29_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_update_completed_
      -- CP-element group 2: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Update/$exit
      -- CP-element group 2: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Update/ack
      -- 
    ack_19_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_29_inst_ack_1, ack => timer_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_sample_completed_
      -- CP-element group 3: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_update_start_
      -- CP-element group 3: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Sample/ra
      -- CP-element group 3: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Update/$entry
      -- CP-element group 3: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Update/cr
      -- 
    ra_28_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_34_inst_ack_0, ack => timer_CP_0_elements(3)); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(3), ack => RPIPE_timer_resp_34_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_update_completed_
      -- CP-element group 4: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Update/$exit
      -- CP-element group 4: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Update/ca
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_34_inst_ack_1, ack => timer_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_32_to_assign_stmt_35/$exit
      -- 
    timer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "timer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timer_CP_0_elements(4) & timer_CP_0_elements(2);
      gj_timer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timer_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal type_cast_31_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_31_wire_constant <= "1";
    -- shared inport operator group (0) : RPIPE_timer_resp_34_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_resp_34_inst_req_0;
      RPIPE_timer_resp_34_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_resp_34_inst_req_1;
      RPIPE_timer_resp_34_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      T_buffer <= data_out(63 downto 0);
      timer_resp_read_0_gI: SplitGuardInterface generic map(name => "timer_resp_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_resp_read_0: InputPortRevised -- 
        generic map ( name => "timer_resp_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_resp_pipe_read_req(0),
          oack => timer_resp_pipe_read_ack(0),
          odata => timer_resp_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_req_29_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_req_29_inst_req_0;
      WPIPE_timer_req_29_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_req_29_inst_req_1;
      WPIPE_timer_req_29_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_31_wire_constant;
      timer_req_write_0_gI: SplitGuardInterface generic map(name => "timer_req_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_req_write_0: OutputPortRevised -- 
        generic map ( name => "timer_req", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_req_pipe_write_req(0),
          oack => timer_req_pipe_write_ack(0),
          odata => timer_req_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_7786_start: Boolean;
  signal timerDaemon_CP_7786_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_2954_branch_req_0 : boolean;
  signal phi_stmt_2956_req_0 : boolean;
  signal phi_stmt_2956_req_1 : boolean;
  signal phi_stmt_2956_ack_0 : boolean;
  signal nCOUNTER_2969_2958_buf_req_0 : boolean;
  signal nCOUNTER_2969_2958_buf_ack_0 : boolean;
  signal nCOUNTER_2969_2958_buf_req_1 : boolean;
  signal nCOUNTER_2969_2958_buf_ack_1 : boolean;
  signal RPIPE_timer_req_2963_inst_req_0 : boolean;
  signal RPIPE_timer_req_2963_inst_ack_0 : boolean;
  signal RPIPE_timer_req_2963_inst_req_1 : boolean;
  signal RPIPE_timer_req_2963_inst_ack_1 : boolean;
  signal WPIPE_timer_resp_2971_inst_req_0 : boolean;
  signal WPIPE_timer_resp_2971_inst_ack_0 : boolean;
  signal WPIPE_timer_resp_2971_inst_req_1 : boolean;
  signal WPIPE_timer_resp_2971_inst_ack_1 : boolean;
  signal do_while_stmt_2954_branch_ack_0 : boolean;
  signal do_while_stmt_2954_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_7786_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_7786_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_7786_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_7786_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_7786: Block -- control-path 
    signal timerDaemon_CP_7786_elements: BooleanArray(44 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_7786_elements(0) <= timerDaemon_CP_7786_start;
    timerDaemon_CP_7786_symbol <= timerDaemon_CP_7786_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2953/$entry
      -- CP-element group 0: 	 branch_block_stmt_2953/branch_block_stmt_2953__entry__
      -- CP-element group 0: 	 branch_block_stmt_2953/do_while_stmt_2954__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	44 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_2953/$exit
      -- CP-element group 1: 	 branch_block_stmt_2953/branch_block_stmt_2953__exit__
      -- CP-element group 1: 	 branch_block_stmt_2953/do_while_stmt_2954__exit__
      -- 
    timerDaemon_CP_7786_elements(1) <= timerDaemon_CP_7786_elements(44);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_2953/do_while_stmt_2954/$entry
      -- CP-element group 2: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954__entry__
      -- 
    timerDaemon_CP_7786_elements(2) <= timerDaemon_CP_7786_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	44 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954__exit__
      -- 
    -- Element group timerDaemon_CP_7786_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_2953/do_while_stmt_2954/loop_back
      -- 
    -- Element group timerDaemon_CP_7786_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	43 
    -- CP-element group 5: 	42 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2953/do_while_stmt_2954/condition_done
      -- CP-element group 5: 	 branch_block_stmt_2953/do_while_stmt_2954/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_2953/do_while_stmt_2954/loop_taken/$entry
      -- 
    timerDaemon_CP_7786_elements(5) <= timerDaemon_CP_7786_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	41 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_2953/do_while_stmt_2954/loop_body_done
      -- 
    timerDaemon_CP_7786_elements(6) <= timerDaemon_CP_7786_elements(41);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_7786_elements(7) <= timerDaemon_CP_7786_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_7786_elements(8) <= timerDaemon_CP_7786_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	40 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/phi_stmt_2961_sample_start_
      -- 
    -- Element group timerDaemon_CP_7786_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	40 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/condition_evaluated
      -- 
    condition_evaluated_7810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_7810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_7786_elements(10), ack => do_while_stmt_2954_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_7786_elements(40) & timerDaemon_CP_7786_elements(14);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7786_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	9 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/phi_stmt_2956_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_7786_elements(15) & timerDaemon_CP_7786_elements(9) & timerDaemon_CP_7786_elements(14);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7786_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	17 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	41 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/phi_stmt_2956_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/phi_stmt_2961_sample_completed_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_7786_elements(35) & timerDaemon_CP_7786_elements(17);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7786_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	32 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/phi_stmt_2956_update_start__ps
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_7786_elements(16) & timerDaemon_CP_7786_elements(32);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7786_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	18 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/aggregated_phi_update_ack
      -- 
    timerDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_7786_elements(36) & timerDaemon_CP_7786_elements(18);
      gj_timerDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7786_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/phi_stmt_2956_sample_start_
      -- 
    timerDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_7786_elements(9) & timerDaemon_CP_7786_elements(12);
      gj_timerDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7786_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	38 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/phi_stmt_2956_update_start_
      -- 
    timerDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_7786_elements(9) & timerDaemon_CP_7786_elements(38);
      gj_timerDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7786_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/phi_stmt_2956_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_7786_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	37 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/phi_stmt_2956_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/phi_stmt_2956_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_7786_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/phi_stmt_2956_loopback_trigger
      -- 
    timerDaemon_CP_7786_elements(19) <= timerDaemon_CP_7786_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/phi_stmt_2956_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/phi_stmt_2956_loopback_sample_req_ps
      -- 
    phi_stmt_2956_loopback_sample_req_7825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2956_loopback_sample_req_7825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_7786_elements(20), ack => phi_stmt_2956_req_0); -- 
    -- Element group timerDaemon_CP_7786_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/phi_stmt_2956_entry_trigger
      -- 
    timerDaemon_CP_7786_elements(21) <= timerDaemon_CP_7786_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/phi_stmt_2956_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/phi_stmt_2956_entry_sample_req_ps
      -- 
    phi_stmt_2956_entry_sample_req_7828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2956_entry_sample_req_7828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_7786_elements(22), ack => phi_stmt_2956_req_1); -- 
    -- Element group timerDaemon_CP_7786_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/phi_stmt_2956_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/phi_stmt_2956_phi_mux_ack_ps
      -- 
    phi_stmt_2956_phi_mux_ack_7831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2956_ack_0, ack => timerDaemon_CP_7786_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/R_nCOUNTER_2958_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/R_nCOUNTER_2958_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/R_nCOUNTER_2958_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/R_nCOUNTER_2958_Sample/req
      -- 
    req_7844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_7786_elements(24), ack => nCOUNTER_2969_2958_buf_req_0); -- 
    -- Element group timerDaemon_CP_7786_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/R_nCOUNTER_2958_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/R_nCOUNTER_2958_update_start_
      -- CP-element group 25: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/R_nCOUNTER_2958_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/R_nCOUNTER_2958_Update/req
      -- 
    req_7849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_7786_elements(25), ack => nCOUNTER_2969_2958_buf_req_1); -- 
    -- Element group timerDaemon_CP_7786_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/R_nCOUNTER_2958_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/R_nCOUNTER_2958_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/R_nCOUNTER_2958_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/R_nCOUNTER_2958_Sample/ack
      -- 
    ack_7845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_2969_2958_buf_ack_0, ack => timerDaemon_CP_7786_elements(26)); -- 
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/R_nCOUNTER_2958_update_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/R_nCOUNTER_2958_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/R_nCOUNTER_2958_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/R_nCOUNTER_2958_Update/ack
      -- 
    ack_7850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_2969_2958_buf_ack_1, ack => timerDaemon_CP_7786_elements(27)); -- 
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/type_cast_2960_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/type_cast_2960_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/type_cast_2960_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/type_cast_2960_sample_completed_
      -- 
    -- Element group timerDaemon_CP_7786_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/type_cast_2960_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/type_cast_2960_update_start_
      -- 
    -- Element group timerDaemon_CP_7786_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/type_cast_2960_update_completed__ps
      -- 
    timerDaemon_CP_7786_elements(30) <= timerDaemon_CP_7786_elements(31);
    -- CP-element group 31:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	30 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/type_cast_2960_update_completed_
      -- 
    -- Element group timerDaemon_CP_7786_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => timerDaemon_CP_7786_elements(29), ack => timerDaemon_CP_7786_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	38 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/phi_stmt_2961_update_start_
      -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_7786_elements(9) & timerDaemon_CP_7786_elements(38);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7786_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/RPIPE_timer_req_2963_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/RPIPE_timer_req_2963_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/RPIPE_timer_req_2963_Sample/rr
      -- 
    rr_7871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_7786_elements(33), ack => RPIPE_timer_req_2963_inst_req_0); -- 
    timerDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_7786_elements(11) & timerDaemon_CP_7786_elements(36);
      gj_timerDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7786_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	13 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/RPIPE_timer_req_2963_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/RPIPE_timer_req_2963_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/RPIPE_timer_req_2963_Update/cr
      -- 
    cr_7876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_7786_elements(34), ack => RPIPE_timer_req_2963_inst_req_1); -- 
    timerDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_7786_elements(35) & timerDaemon_CP_7786_elements(13);
      gj_timerDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7786_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/RPIPE_timer_req_2963_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/RPIPE_timer_req_2963_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/RPIPE_timer_req_2963_Sample/ra
      -- 
    ra_7872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_2963_inst_ack_0, ack => timerDaemon_CP_7786_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	37 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/phi_stmt_2961_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/RPIPE_timer_req_2963_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/RPIPE_timer_req_2963_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/RPIPE_timer_req_2963_Update/ca
      -- 
    ca_7877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_2963_inst_ack_1, ack => timerDaemon_CP_7786_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: 	18 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/WPIPE_timer_resp_2971_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/WPIPE_timer_resp_2971_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/WPIPE_timer_resp_2971_Sample/req
      -- 
    req_7885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_7786_elements(37), ack => WPIPE_timer_resp_2971_inst_req_0); -- 
    timerDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_7786_elements(36) & timerDaemon_CP_7786_elements(18) & timerDaemon_CP_7786_elements(39);
      gj_timerDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7786_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	16 
    -- CP-element group 38: 	32 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/WPIPE_timer_resp_2971_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/WPIPE_timer_resp_2971_update_start_
      -- CP-element group 38: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/WPIPE_timer_resp_2971_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/WPIPE_timer_resp_2971_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/WPIPE_timer_resp_2971_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/WPIPE_timer_resp_2971_Update/req
      -- 
    ack_7886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_2971_inst_ack_0, ack => timerDaemon_CP_7786_elements(38)); -- 
    req_7890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_7786_elements(38), ack => WPIPE_timer_resp_2971_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/WPIPE_timer_resp_2971_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/WPIPE_timer_resp_2971_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/WPIPE_timer_resp_2971_Update/ack
      -- 
    ack_7891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_2971_inst_ack_1, ack => timerDaemon_CP_7786_elements(39)); -- 
    -- CP-element group 40:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	10 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_7786_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => timerDaemon_CP_7786_elements(9), ack => timerDaemon_CP_7786_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: 	12 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	6 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_2953/do_while_stmt_2954/do_while_stmt_2954_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_7786_elements(39) & timerDaemon_CP_7786_elements(12);
      gj_timerDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7786_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	5 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_2953/do_while_stmt_2954/loop_exit/$exit
      -- CP-element group 42: 	 branch_block_stmt_2953/do_while_stmt_2954/loop_exit/ack
      -- 
    ack_7896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2954_branch_ack_0, ack => timerDaemon_CP_7786_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	5 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_2953/do_while_stmt_2954/loop_taken/$exit
      -- CP-element group 43: 	 branch_block_stmt_2953/do_while_stmt_2954/loop_taken/ack
      -- 
    ack_7900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2954_branch_ack_1, ack => timerDaemon_CP_7786_elements(43)); -- 
    -- CP-element group 44:  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	3 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	1 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_2953/do_while_stmt_2954/$exit
      -- 
    timerDaemon_CP_7786_elements(44) <= timerDaemon_CP_7786_elements(3);
    timerDaemon_do_while_stmt_2954_terminator_7901: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_2954_terminator_7901", max_iterations_in_flight =>7) 
      port map(loop_body_exit => timerDaemon_CP_7786_elements(6),loop_continue => timerDaemon_CP_7786_elements(43),loop_terminate => timerDaemon_CP_7786_elements(42),loop_back => timerDaemon_CP_7786_elements(4),loop_exit => timerDaemon_CP_7786_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_2956_phi_seq_7859_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_7786_elements(19);
      timerDaemon_CP_7786_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_7786_elements(26);
      timerDaemon_CP_7786_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_7786_elements(27);
      timerDaemon_CP_7786_elements(20) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_7786_elements(21);
      timerDaemon_CP_7786_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_7786_elements(28);
      timerDaemon_CP_7786_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_7786_elements(30);
      timerDaemon_CP_7786_elements(22) <= phi_mux_reqs(1);
      phi_stmt_2956_phi_seq_7859 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_2956_phi_seq_7859") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_7786_elements(11), 
          phi_sample_ack => timerDaemon_CP_7786_elements(17), 
          phi_update_req => timerDaemon_CP_7786_elements(13), 
          phi_update_ack => timerDaemon_CP_7786_elements(18), 
          phi_mux_ack => timerDaemon_CP_7786_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_7811_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_7786_elements(7);
        preds(1)  <= timerDaemon_CP_7786_elements(8);
        entry_tmerge_7811 : transition_merge -- 
          generic map(name => " entry_tmerge_7811")
          port map (preds => preds, symbol_out => timerDaemon_CP_7786_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal COUNTER_2956 : std_logic_vector(63 downto 0);
    signal RPIPE_timer_req_2963_wire : std_logic_vector(0 downto 0);
    signal konst_2967_wire_constant : std_logic_vector(63 downto 0);
    signal konst_2975_wire_constant : std_logic_vector(0 downto 0);
    signal nCOUNTER_2969 : std_logic_vector(63 downto 0);
    signal nCOUNTER_2969_2958_buffered : std_logic_vector(63 downto 0);
    signal req_2961 : std_logic_vector(0 downto 0);
    signal type_cast_2960_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_2967_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_2975_wire_constant <= "1";
    type_cast_2960_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_2956: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nCOUNTER_2969_2958_buffered & type_cast_2960_wire_constant;
      req <= phi_stmt_2956_req_0 & phi_stmt_2956_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2956",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2956_ack_0,
          idata => idata,
          odata => COUNTER_2956,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2956
    nCOUNTER_2969_2958_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nCOUNTER_2969_2958_buf_req_0;
      nCOUNTER_2969_2958_buf_ack_0<= wack(0);
      rreq(0) <= nCOUNTER_2969_2958_buf_req_1;
      nCOUNTER_2969_2958_buf_ack_1<= rack(0);
      nCOUNTER_2969_2958_buf : InterlockBuffer generic map ( -- 
        name => "nCOUNTER_2969_2958_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nCOUNTER_2969,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nCOUNTER_2969_2958_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_2961
    process(RPIPE_timer_req_2963_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := RPIPE_timer_req_2963_wire(0 downto 0);
      req_2961 <= tmp_var; -- 
    end process;
    do_while_stmt_2954_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_2975_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2954_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2954_branch_req_0,
          ack0 => do_while_stmt_2954_branch_ack_0,
          ack1 => do_while_stmt_2954_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_2968_inst
    process(COUNTER_2956) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(COUNTER_2956, konst_2967_wire_constant, tmp_var);
      nCOUNTER_2969 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_timer_req_2963_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_req_2963_inst_req_0;
      RPIPE_timer_req_2963_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_req_2963_inst_req_1;
      RPIPE_timer_req_2963_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_timer_req_2963_wire <= data_out(0 downto 0);
      timer_req_read_0_gI: SplitGuardInterface generic map(name => "timer_req_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_req_read_0: InputPortRevised -- 
        generic map ( name => "timer_req_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_req_pipe_read_req(0),
          oack => timer_req_pipe_read_ack(0),
          odata => timer_req_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_resp_2971_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_resp_2971_inst_req_0;
      WPIPE_timer_resp_2971_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_resp_2971_inst_req_1;
      WPIPE_timer_resp_2971_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= req_2961(0);
      data_in <= COUNTER_2956;
      timer_resp_write_0_gI: SplitGuardInterface generic map(name => "timer_resp_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_resp_write_0: OutputPortRevised -- 
        generic map ( name => "timer_resp", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_resp_pipe_write_req(0),
          oack => timer_resp_pipe_write_ack(0),
          odata => timer_resp_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(69 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(319 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(94 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(4 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_T :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_start
  signal Block2_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_start
  signal Block3_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_req
  signal timer_req_pipe_write_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_req
  signal timer_req_pipe_read_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_resp
  signal timer_resp_pipe_write_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_resp
  signal timer_resp_pipe_read_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(18 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(18 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(10 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(0 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(4 downto 4),
      memory_space_2_sr_ack => memory_space_2_sr_ack(4 downto 4),
      memory_space_2_sr_addr => memory_space_2_sr_addr(69 downto 56),
      memory_space_2_sr_data => memory_space_2_sr_data(319 downto 256),
      memory_space_2_sr_tag => memory_space_2_sr_tag(94 downto 76),
      memory_space_2_sc_req => memory_space_2_sc_req(4 downto 4),
      memory_space_2_sc_ack => memory_space_2_sc_ack(4 downto 4),
      memory_space_2_sc_tag => memory_space_2_sc_tag(4 downto 4),
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(15 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(15 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(15 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(15 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(15 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(15 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(3 downto 3),
      memory_space_0_lr_ack => memory_space_0_lr_ack(3 downto 3),
      memory_space_0_lr_addr => memory_space_0_lr_addr(55 downto 42),
      memory_space_0_lr_tag => memory_space_0_lr_tag(75 downto 57),
      memory_space_0_lc_req => memory_space_0_lc_req(3 downto 3),
      memory_space_0_lc_ack => memory_space_0_lc_ack(3 downto 3),
      memory_space_0_lc_data => memory_space_0_lc_data(255 downto 192),
      memory_space_0_lc_tag => memory_space_0_lc_tag(3 downto 3),
      memory_space_2_sr_req => memory_space_2_sr_req(3 downto 3),
      memory_space_2_sr_ack => memory_space_2_sr_ack(3 downto 3),
      memory_space_2_sr_addr => memory_space_2_sr_addr(55 downto 42),
      memory_space_2_sr_data => memory_space_2_sr_data(255 downto 192),
      memory_space_2_sr_tag => memory_space_2_sr_tag(75 downto 57),
      memory_space_2_sc_req => memory_space_2_sc_req(3 downto 3),
      memory_space_2_sc_ack => memory_space_2_sc_ack(3 downto 3),
      memory_space_2_sc_tag => memory_space_2_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(2 downto 2),
      memory_space_0_lr_ack => memory_space_0_lr_ack(2 downto 2),
      memory_space_0_lr_addr => memory_space_0_lr_addr(41 downto 28),
      memory_space_0_lr_tag => memory_space_0_lr_tag(56 downto 38),
      memory_space_0_lc_req => memory_space_0_lc_req(2 downto 2),
      memory_space_0_lc_ack => memory_space_0_lc_ack(2 downto 2),
      memory_space_0_lc_data => memory_space_0_lc_data(191 downto 128),
      memory_space_0_lc_tag => memory_space_0_lc_tag(2 downto 2),
      memory_space_2_sr_req => memory_space_2_sr_req(2 downto 2),
      memory_space_2_sr_ack => memory_space_2_sr_ack(2 downto 2),
      memory_space_2_sr_addr => memory_space_2_sr_addr(41 downto 28),
      memory_space_2_sr_data => memory_space_2_sr_data(191 downto 128),
      memory_space_2_sr_tag => memory_space_2_sr_tag(56 downto 38),
      memory_space_2_sc_req => memory_space_2_sc_req(2 downto 2),
      memory_space_2_sc_ack => memory_space_2_sc_ack(2 downto 2),
      memory_space_2_sc_tag => memory_space_2_sc_tag(2 downto 2),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(15 downto 0),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(18 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(13 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(18 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      Block2_start_pipe_read_req => Block2_start_pipe_read_req(0 downto 0),
      Block2_start_pipe_read_ack => Block2_start_pipe_read_ack(0 downto 0),
      Block2_start_pipe_read_data => Block2_start_pipe_read_data(15 downto 0),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(27 downto 14),
      memory_space_0_lr_tag => memory_space_0_lr_tag(37 downto 19),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(127 downto 64),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 1),
      memory_space_2_sr_req => memory_space_2_sr_req(1 downto 1),
      memory_space_2_sr_ack => memory_space_2_sr_ack(1 downto 1),
      memory_space_2_sr_addr => memory_space_2_sr_addr(27 downto 14),
      memory_space_2_sr_data => memory_space_2_sr_data(127 downto 64),
      memory_space_2_sr_tag => memory_space_2_sr_tag(37 downto 19),
      memory_space_2_sc_req => memory_space_2_sc_req(1 downto 1),
      memory_space_2_sc_ack => memory_space_2_sc_ack(1 downto 1),
      memory_space_2_sc_tag => memory_space_2_sc_tag(1 downto 1),
      Block3_start_pipe_read_req => Block3_start_pipe_read_req(0 downto 0),
      Block3_start_pipe_read_ack => Block3_start_pipe_read_ack(0 downto 0),
      Block3_start_pipe_read_data => Block3_start_pipe_read_data(15 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module timer
  timer_out_args <= timer_T ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      T => timer_T,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      timer_resp_pipe_read_req => timer_resp_pipe_read_req(0 downto 0),
      timer_resp_pipe_read_ack => timer_resp_pipe_read_ack(0 downto 0),
      timer_resp_pipe_read_data => timer_resp_pipe_read_data(63 downto 0),
      timer_req_pipe_write_req => timer_req_pipe_write_req(0 downto 0),
      timer_req_pipe_write_ack => timer_req_pipe_write_ack(0 downto 0),
      timer_req_pipe_write_data => timer_req_pipe_write_data(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      timer_req_pipe_read_req => timer_req_pipe_read_req(0 downto 0),
      timer_req_pipe_read_ack => timer_req_pipe_read_ack(0 downto 0),
      timer_req_pipe_read_data => timer_req_pipe_read_data(0 downto 0),
      timer_resp_pipe_write_req => timer_resp_pipe_write_req(0 downto 0),
      timer_resp_pipe_write_ack => timer_resp_pipe_write_ack(0 downto 0),
      timer_resp_pipe_write_data => timer_resp_pipe_write_data(63 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  timer_req_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_req",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_req_pipe_read_req,
      read_ack => timer_req_pipe_read_ack,
      read_data => timer_req_pipe_read_data,
      write_req => timer_req_pipe_write_req,
      write_ack => timer_req_pipe_write_ack,
      write_data => timer_req_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  timer_resp_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_resp",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_resp_pipe_read_req,
      read_ack => timer_resp_pipe_read_ack,
      read_data => timer_resp_pipe_read_data,
      write_req => timer_resp_pipe_write_req,
      write_ack => timer_resp_pipe_write_ack,
      write_data => timer_resp_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_1: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 5,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
